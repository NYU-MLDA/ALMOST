//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n955_, new_n957_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_;
  XOR2_X1   g000(.A(G71gat), .B(G99gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT81), .B(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G15gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n204_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT25), .B(G183gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(KEYINPUT24), .A3(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n211_), .A2(new_n216_), .A3(new_n220_), .A4(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n214_), .B(new_n215_), .C1(G183gat), .C2(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n221_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT79), .B(G176gat), .Z(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT22), .B(G169gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n224_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  AOI211_X1 g029(.A(KEYINPUT80), .B(new_n225_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n223_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT30), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n208_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n208_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n240_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  OR3_X1    g048(.A1(new_n237_), .A2(new_n239_), .A3(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT27), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT19), .ZN(new_n255_));
  INV_X1    g054(.A(G197gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G204gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT21), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(KEYINPUT86), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT85), .B(G204gat), .Z(new_n260_));
  OAI211_X1 g059(.A(new_n257_), .B(new_n259_), .C1(new_n260_), .C2(new_n256_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G211gat), .B(G218gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(G204gat), .B1(new_n256_), .B2(KEYINPUT86), .ZN(new_n263_));
  NAND2_X1  g062(.A1(KEYINPUT86), .A2(G197gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n261_), .B(new_n262_), .C1(new_n265_), .C2(new_n258_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT87), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n257_), .B1(new_n260_), .B2(new_n256_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n262_), .A2(new_n258_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n266_), .A2(new_n267_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n267_), .B1(new_n266_), .B2(new_n270_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n271_), .A2(new_n272_), .A3(new_n232_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n226_), .A2(new_n227_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT89), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n221_), .B(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n224_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT90), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n274_), .A2(new_n224_), .A3(KEYINPUT90), .A4(new_n276_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n223_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n266_), .A2(new_n270_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT20), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n255_), .B1(new_n273_), .B2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286_));
  INV_X1    g085(.A(G92gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT18), .B(G64gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n232_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n281_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n282_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT91), .B1(new_n281_), .B2(new_n282_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n255_), .A2(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n291_), .A2(new_n295_), .A3(new_n296_), .A4(new_n298_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n285_), .A2(new_n290_), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n290_), .B1(new_n285_), .B2(new_n299_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n253_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n297_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n282_), .A2(KEYINPUT87), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n266_), .A2(new_n267_), .A3(new_n270_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n303_), .B1(new_n306_), .B2(new_n232_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n255_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n297_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n277_), .A2(new_n223_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT95), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n314_), .B2(new_n293_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n291_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n290_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n309_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n285_), .A2(new_n299_), .A3(new_n290_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT27), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n302_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT92), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324_));
  INV_X1    g123(.A(G141gat), .ZN(new_n325_));
  INV_X1    g124(.A(G148gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT2), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n327_), .A2(new_n330_), .A3(new_n331_), .A4(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(KEYINPUT1), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G155gat), .A3(G162gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n340_), .A3(new_n334_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G141gat), .B(G148gat), .Z(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n323_), .B1(new_n344_), .B2(new_n246_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n243_), .A2(new_n245_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n333_), .A2(new_n336_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(new_n323_), .A3(new_n347_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n322_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n346_), .A2(new_n347_), .A3(KEYINPUT4), .ZN(new_n353_));
  OR3_X1    g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G1gat), .B(G29gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT93), .B(G85gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT0), .B(G57gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n352_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n354_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n359_), .B1(new_n365_), .B2(new_n362_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G78gat), .B(G106gat), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n344_), .A2(KEYINPUT29), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G228gat), .A2(G233gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n371_), .B1(new_n282_), .B2(new_n370_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n369_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  OR3_X1    g174(.A1(new_n344_), .A2(KEYINPUT84), .A3(KEYINPUT29), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT84), .B1(new_n344_), .B2(KEYINPUT29), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G22gat), .B(G50gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT28), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n372_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n282_), .A2(new_n370_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n371_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n368_), .A3(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n375_), .A2(new_n382_), .A3(KEYINPUT88), .A4(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT88), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n392_), .A2(new_n382_), .B1(new_n388_), .B2(new_n375_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  NOR4_X1   g193(.A1(new_n252_), .A2(new_n321_), .A3(new_n367_), .A4(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n367_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT96), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n302_), .A4(new_n320_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(new_n382_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n375_), .A2(new_n388_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n401_), .A2(new_n366_), .A3(new_n364_), .A4(new_n389_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT96), .B1(new_n321_), .B2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n365_), .A2(new_n362_), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT33), .B1(new_n404_), .B2(new_n360_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  NOR4_X1   g205(.A1(new_n365_), .A2(new_n406_), .A3(new_n359_), .A4(new_n362_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n349_), .A2(new_n350_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n359_), .B1(new_n410_), .B2(new_n352_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n351_), .A2(new_n361_), .A3(new_n353_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n300_), .A2(new_n301_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n290_), .A2(KEYINPUT32), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n285_), .A2(new_n299_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT94), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT94), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n285_), .A2(new_n299_), .A3(new_n418_), .A4(new_n415_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n307_), .A2(new_n308_), .B1(new_n315_), .B2(new_n291_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n415_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n364_), .A2(new_n366_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n408_), .A2(new_n414_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n398_), .B(new_n403_), .C1(new_n394_), .C2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n395_), .B1(new_n425_), .B2(new_n252_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT13), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT65), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G85gat), .A2(G92gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT64), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n430_), .B1(new_n431_), .B2(KEYINPUT9), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT9), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(KEYINPUT64), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n429_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n430_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G85gat), .A2(G92gat), .ZN(new_n437_));
  OAI22_X1  g236(.A1(new_n436_), .A2(new_n437_), .B1(KEYINPUT9), .B2(new_n287_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n431_), .A2(KEYINPUT9), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(KEYINPUT64), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT65), .A4(new_n430_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n435_), .A2(new_n438_), .A3(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(KEYINPUT10), .B(G99gat), .Z(new_n443_));
  INV_X1    g242(.A(G106gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G99gat), .A2(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT6), .ZN(new_n446_));
  AND2_X1   g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n443_), .A2(new_n444_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n442_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT8), .ZN(new_n452_));
  AND2_X1   g251(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n453_));
  NOR2_X1   g252(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n445_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT66), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n448_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n447_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n460_));
  OR3_X1    g259(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n455_), .A2(new_n459_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n436_), .A2(new_n437_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n452_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n452_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n461_), .A2(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n449_), .A2(new_n446_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n451_), .B1(new_n464_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G57gat), .ZN(new_n470_));
  INV_X1    g269(.A(G64gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G57gat), .A2(G64gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT11), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G71gat), .B(G78gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT11), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n472_), .A2(new_n478_), .A3(new_n473_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n475_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n476_), .A3(KEYINPUT11), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n469_), .A2(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n451_), .B(new_n482_), .C1(new_n464_), .C2(new_n468_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G230gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n485_), .A2(KEYINPUT67), .A3(new_n487_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT67), .B1(new_n485_), .B2(new_n487_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT12), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n484_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n469_), .A2(KEYINPUT12), .A3(new_n483_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n492_), .A2(new_n496_), .A3(KEYINPUT68), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT68), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n485_), .A2(new_n487_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n485_), .A2(KEYINPUT67), .A3(new_n487_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n469_), .A2(KEYINPUT12), .A3(new_n483_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT12), .B1(new_n469_), .B2(new_n483_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n498_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n489_), .B1(new_n497_), .B2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n509_));
  XNOR2_X1  g308(.A(G120gat), .B(G148gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G176gat), .B(G204gat), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n511_), .B(new_n512_), .Z(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n513_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n489_), .B(new_n516_), .C1(new_n497_), .C2(new_n507_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n428_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(KEYINPUT13), .A3(new_n517_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT15), .ZN(new_n522_));
  INV_X1    g321(.A(G50gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(G43gat), .ZN(new_n524_));
  INV_X1    g323(.A(G43gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(G50gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n524_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G29gat), .B(G36gat), .Z(new_n530_));
  NOR3_X1   g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G29gat), .B(G36gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n525_), .A2(G50gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n523_), .A2(G43gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT70), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n524_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n532_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n522_), .B1(new_n531_), .B2(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(G1gat), .A2(G8gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G1gat), .A2(G8gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(G15gat), .A2(G22gat), .ZN(new_n542_));
  NOR2_X1   g341(.A1(G15gat), .A2(G22gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(G1gat), .B2(G8gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n541_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n548_), .A2(new_n545_), .A3(new_n540_), .A4(new_n539_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n530_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n535_), .A2(new_n536_), .A3(new_n532_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT15), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n538_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n550_), .B1(new_n552_), .B2(new_n551_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT77), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT77), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n554_), .A2(new_n556_), .A3(new_n560_), .A4(new_n557_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n551_), .A2(new_n552_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n550_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n562_), .B1(new_n565_), .B2(new_n555_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT76), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(KEYINPUT76), .B(new_n562_), .C1(new_n565_), .C2(new_n555_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n559_), .A2(new_n561_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G169gat), .B(G197gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT78), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n559_), .A2(new_n561_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n568_), .A2(new_n569_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n573_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(KEYINPUT78), .A3(new_n573_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n521_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT73), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT36), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT71), .ZN(new_n593_));
  INV_X1    g392(.A(new_n563_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n469_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n593_), .B1(new_n469_), .B2(new_n594_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n469_), .A2(new_n553_), .A3(new_n538_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT34), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT35), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .A4(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n600_), .A2(new_n601_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT72), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(new_n606_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n603_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n608_), .B1(new_n603_), .B2(new_n609_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n592_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n590_), .B(KEYINPUT36), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n610_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT37), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n613_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n615_), .B(KEYINPUT74), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(new_n610_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n617_), .B1(new_n613_), .B2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n550_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(new_n482_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G127gat), .B(G155gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(G211gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT16), .B(G183gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(KEYINPUT17), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n625_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(KEYINPUT17), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n625_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(KEYINPUT75), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(KEYINPUT75), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n622_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n427_), .A2(new_n586_), .A3(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n364_), .A2(new_n366_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n640_), .A2(G1gat), .A3(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT97), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n643_), .A2(KEYINPUT38), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(KEYINPUT38), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n613_), .A2(new_n616_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT98), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT98), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(new_n637_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n427_), .A2(new_n586_), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n641_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n644_), .A2(new_n645_), .A3(new_n652_), .ZN(G1324gat));
  INV_X1    g452(.A(new_n321_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT99), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n658_), .B(G8gat), .C1(new_n651_), .C2(new_n654_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(KEYINPUT39), .A3(new_n659_), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n640_), .A2(G8gat), .A3(new_n654_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT39), .B1(new_n657_), .B2(new_n659_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n665_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n662_), .A2(new_n663_), .A3(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1325gat));
  OAI21_X1  g468(.A(G15gat), .B1(new_n651_), .B2(new_n252_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n670_), .A2(KEYINPUT41), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(KEYINPUT41), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n640_), .A2(G15gat), .A3(new_n252_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n671_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT101), .Z(G1326gat));
  INV_X1    g474(.A(new_n394_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G22gat), .B1(new_n651_), .B2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n678_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n676_), .A2(G22gat), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT103), .Z(new_n682_));
  OAI211_X1 g481(.A(new_n679_), .B(new_n680_), .C1(new_n640_), .C2(new_n682_), .ZN(G1327gat));
  NOR2_X1   g482(.A1(new_n646_), .A2(new_n637_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n252_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n417_), .A2(new_n419_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n421_), .A2(new_n422_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n367_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n364_), .A2(new_n406_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n404_), .A2(KEYINPUT33), .A3(new_n360_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n285_), .A2(new_n299_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n317_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n413_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n319_), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n686_), .A2(new_n688_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n394_), .A2(new_n302_), .A3(new_n320_), .A4(new_n641_), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n696_), .A2(new_n676_), .B1(new_n697_), .B2(KEYINPUT96), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n685_), .B1(new_n698_), .B2(new_n398_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n586_), .B(new_n684_), .C1(new_n699_), .C2(new_n395_), .ZN(new_n700_));
  OR3_X1    g499(.A1(new_n700_), .A2(G29gat), .A3(new_n641_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n622_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n426_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n704_), .B(new_n622_), .C1(new_n699_), .C2(new_n395_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n586_), .A3(new_n638_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n637_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(KEYINPUT44), .A3(new_n586_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(new_n367_), .A3(new_n711_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n712_), .A2(KEYINPUT104), .A3(G29gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT104), .B1(new_n712_), .B2(G29gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n701_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  NAND3_X1  g514(.A1(new_n709_), .A2(new_n321_), .A3(new_n711_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G36gat), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719_));
  INV_X1    g518(.A(new_n521_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n584_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n684_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n426_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n654_), .A2(G36gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n719_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n724_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n700_), .A2(KEYINPUT105), .A3(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n718_), .B1(new_n725_), .B2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n723_), .A2(new_n719_), .A3(new_n724_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT105), .B1(new_n700_), .B2(new_n726_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(KEYINPUT45), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n717_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT46), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n732_), .B1(new_n716_), .B2(G36gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n737_), .A2(KEYINPUT106), .A3(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1329gat));
  NAND4_X1  g539(.A1(new_n709_), .A2(G43gat), .A3(new_n685_), .A4(new_n711_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G43gat), .B1(new_n723_), .B2(new_n685_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT107), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g544(.A1(new_n723_), .A2(new_n523_), .A3(new_n394_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n709_), .A2(new_n394_), .A3(new_n711_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(new_n523_), .ZN(G1331gat));
  NOR2_X1   g547(.A1(new_n720_), .A2(new_n584_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(new_n426_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n650_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n752_), .A2(new_n470_), .A3(new_n641_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(KEYINPUT108), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(KEYINPUT108), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n751_), .A2(new_n639_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G57gat), .B1(new_n758_), .B2(new_n367_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n755_), .A2(new_n756_), .A3(new_n759_), .ZN(G1332gat));
  OAI21_X1  g559(.A(G64gat), .B1(new_n752_), .B2(new_n654_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT48), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(new_n471_), .A3(new_n321_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1333gat));
  OAI21_X1  g563(.A(G71gat), .B1(new_n752_), .B2(new_n252_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT49), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n252_), .A2(G71gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n757_), .B2(new_n767_), .ZN(G1334gat));
  OAI21_X1  g567(.A(G78gat), .B1(new_n752_), .B2(new_n676_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT50), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n676_), .A2(G78gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n757_), .B2(new_n771_), .ZN(G1335gat));
  NOR3_X1   g571(.A1(new_n750_), .A2(new_n426_), .A3(new_n722_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n367_), .ZN(new_n774_));
  INV_X1    g573(.A(G85gat), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT109), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n706_), .A2(KEYINPUT110), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n703_), .A2(new_n705_), .A3(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n750_), .A2(new_n637_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n778_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(G85gat), .A3(new_n367_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n777_), .A2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT111), .ZN(G1336gat));
  AOI21_X1  g584(.A(G92gat), .B1(new_n773_), .B2(new_n321_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n654_), .A2(new_n287_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n782_), .B2(new_n787_), .ZN(G1337gat));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n789_), .A2(KEYINPUT112), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n778_), .A2(new_n685_), .A3(new_n780_), .A4(new_n781_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G99gat), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n685_), .A2(new_n443_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n773_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n790_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n794_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n789_), .A2(KEYINPUT113), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n790_), .B2(KEYINPUT113), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n796_), .B(new_n798_), .C1(new_n791_), .C2(G99gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT114), .B1(new_n795_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n798_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n792_), .A2(new_n794_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n796_), .B1(new_n791_), .B2(G99gat), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n802_), .B(new_n803_), .C1(new_n804_), .C2(new_n790_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n800_), .A2(new_n805_), .ZN(G1338gat));
  NAND3_X1  g605(.A1(new_n773_), .A2(new_n444_), .A3(new_n394_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n750_), .A2(new_n676_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n710_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n810_), .B2(G106gat), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT52), .B(new_n444_), .C1(new_n710_), .C2(new_n809_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n807_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g613(.A1(new_n252_), .A2(new_n394_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n321_), .A2(new_n641_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n570_), .A2(new_n574_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n554_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n565_), .A2(new_n555_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n820_), .B(new_n573_), .C1(new_n821_), .C2(new_n562_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n517_), .A2(new_n819_), .A3(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT68), .B1(new_n492_), .B2(new_n496_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n503_), .A2(new_n506_), .A3(new_n498_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT55), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n485_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n488_), .B1(new_n496_), .B2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n503_), .A2(new_n506_), .A3(KEYINPUT55), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n513_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT56), .B(new_n513_), .C1(new_n826_), .C2(new_n830_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n823_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n622_), .B1(new_n835_), .B2(KEYINPUT58), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT117), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n622_), .B(new_n838_), .C1(new_n835_), .C2(KEYINPUT58), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n840_), .B(new_n823_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n837_), .A2(new_n839_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n833_), .A2(new_n834_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n580_), .A2(new_n517_), .A3(new_n582_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n580_), .A2(new_n517_), .A3(KEYINPUT116), .A4(new_n582_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n845_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n819_), .A2(new_n822_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n844_), .B1(new_n854_), .B2(new_n646_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n646_), .ZN(new_n856_));
  AOI211_X1 g655(.A(KEYINPUT57), .B(new_n856_), .C1(new_n850_), .C2(new_n853_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n843_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT118), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n843_), .B(new_n860_), .C1(new_n855_), .C2(new_n857_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n638_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n585_), .A2(new_n637_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n863_), .A2(KEYINPUT115), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n622_), .B1(new_n863_), .B2(KEYINPUT115), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n720_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT54), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n864_), .A2(new_n865_), .A3(new_n868_), .A4(new_n720_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  AOI211_X1 g669(.A(new_n816_), .B(new_n818_), .C1(new_n862_), .C2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(G113gat), .B1(new_n871_), .B2(new_n584_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n818_), .A2(KEYINPUT59), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n858_), .A2(new_n638_), .ZN(new_n875_));
  AOI211_X1 g674(.A(new_n816_), .B(new_n874_), .C1(new_n875_), .C2(new_n870_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n848_), .A2(new_n849_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n852_), .B1(new_n877_), .B2(new_n845_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT57), .B1(new_n878_), .B2(new_n856_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n854_), .A2(new_n844_), .A3(new_n646_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n841_), .B1(new_n836_), .B2(KEYINPUT117), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n879_), .A2(new_n880_), .B1(new_n881_), .B2(new_n839_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n638_), .B1(new_n882_), .B2(new_n860_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n861_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n870_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n876_), .B1(new_n886_), .B2(KEYINPUT59), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n584_), .A2(G113gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n872_), .B1(new_n887_), .B2(new_n888_), .ZN(G1340gat));
  INV_X1    g688(.A(G120gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n720_), .B2(KEYINPUT60), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n871_), .B(new_n891_), .C1(KEYINPUT60), .C2(new_n890_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n720_), .B(new_n876_), .C1(new_n886_), .C2(KEYINPUT59), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n890_), .ZN(G1341gat));
  NAND4_X1  g693(.A1(new_n885_), .A2(new_n815_), .A3(new_n637_), .A4(new_n817_), .ZN(new_n895_));
  INV_X1    g694(.A(G127gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n876_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n638_), .A2(new_n896_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n900_), .B(new_n901_), .C1(new_n871_), .C2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n895_), .A2(KEYINPUT119), .A3(new_n896_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n899_), .A2(new_n903_), .A3(new_n904_), .ZN(G1342gat));
  NAND2_X1  g704(.A1(new_n647_), .A2(new_n648_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G134gat), .B1(new_n871_), .B2(new_n906_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n622_), .A2(G134gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n887_), .B2(new_n908_), .ZN(G1343gat));
  INV_X1    g708(.A(new_n870_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n637_), .B1(new_n858_), .B2(KEYINPUT118), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n861_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n685_), .A2(new_n676_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n817_), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT120), .Z(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n912_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n584_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n521_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT121), .B(G148gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1345gat));
  XNOR2_X1  g721(.A(KEYINPUT61), .B(G155gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n917_), .B2(new_n637_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n885_), .A2(new_n637_), .A3(new_n915_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(KEYINPUT122), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n924_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n917_), .A2(new_n925_), .A3(new_n637_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n927_), .A2(KEYINPUT122), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n930_), .A2(new_n931_), .A3(new_n923_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n929_), .A2(new_n932_), .ZN(G1346gat));
  AND3_X1   g732(.A1(new_n917_), .A2(G162gat), .A3(new_n622_), .ZN(new_n934_));
  AOI21_X1  g733(.A(G162gat), .B1(new_n917_), .B2(new_n906_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1347gat));
  AOI21_X1  g735(.A(new_n816_), .B1(new_n875_), .B2(new_n870_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n654_), .A2(new_n367_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n937_), .A2(new_n584_), .A3(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n939_), .A2(new_n940_), .A3(G169gat), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n939_), .A2(G169gat), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(KEYINPUT62), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n939_), .A2(KEYINPUT123), .A3(new_n940_), .A4(G169gat), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n943_), .A2(new_n945_), .A3(new_n946_), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n937_), .A2(new_n584_), .A3(new_n227_), .A4(new_n938_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1348gat));
  NOR2_X1   g748(.A1(new_n912_), .A2(new_n816_), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n950_), .A2(G176gat), .A3(new_n521_), .A4(new_n938_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n937_), .A2(new_n938_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n226_), .B1(new_n952_), .B2(new_n720_), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1349gat));
  NOR2_X1   g753(.A1(new_n952_), .A2(new_n638_), .ZN(new_n955_));
  MUX2_X1   g754(.A(G183gat), .B(new_n209_), .S(new_n955_), .Z(G1350gat));
  OAI21_X1  g755(.A(G190gat), .B1(new_n952_), .B2(new_n702_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n906_), .A2(new_n210_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(KEYINPUT124), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n957_), .B1(new_n952_), .B2(new_n959_), .ZN(G1351gat));
  NAND2_X1  g759(.A1(new_n913_), .A2(new_n938_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n912_), .A2(new_n961_), .ZN(new_n962_));
  AOI22_X1  g761(.A1(new_n962_), .A2(new_n584_), .B1(KEYINPUT125), .B2(G197gat), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n963_), .B1(KEYINPUT125), .B2(G197gat), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965_));
  NAND4_X1  g764(.A1(new_n962_), .A2(new_n965_), .A3(new_n256_), .A4(new_n584_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n964_), .A2(new_n966_), .ZN(G1352gat));
  OR4_X1    g766(.A1(new_n720_), .A2(new_n912_), .A3(new_n260_), .A4(new_n961_), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n912_), .A2(new_n720_), .A3(new_n961_), .ZN(new_n969_));
  INV_X1    g768(.A(G204gat), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n968_), .B1(new_n969_), .B2(new_n970_), .ZN(G1353gat));
  AOI21_X1  g770(.A(new_n638_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n962_), .A2(new_n972_), .ZN(new_n973_));
  XOR2_X1   g772(.A(KEYINPUT126), .B(KEYINPUT127), .Z(new_n974_));
  NOR2_X1   g773(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n974_), .B(new_n975_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n973_), .B(new_n976_), .ZN(G1354gat));
  AOI21_X1  g776(.A(G218gat), .B1(new_n962_), .B2(new_n906_), .ZN(new_n978_));
  AND2_X1   g777(.A1(new_n622_), .A2(G218gat), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n978_), .B1(new_n962_), .B2(new_n979_), .ZN(G1355gat));
endmodule


