//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n204_), .A2(new_n205_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(KEYINPUT64), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(KEYINPUT64), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n210_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  OAI22_X1  g021(.A1(new_n222_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n205_), .A4(KEYINPUT65), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n208_), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n223_), .B(new_n226_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n215_), .A2(new_n218_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n221_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G57gat), .B(G64gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G78gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n239_));
  XOR2_X1   g038(.A(G71gat), .B(G78gat), .Z(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(KEYINPUT11), .A3(new_n235_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n238_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n234_), .A2(new_n243_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n242_), .B(new_n221_), .C1(new_n233_), .C2(new_n232_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT12), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT12), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n234_), .A2(new_n247_), .A3(new_n243_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n203_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n202_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G120gat), .B(G148gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT5), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G176gat), .ZN(new_n254_));
  INV_X1    g053(.A(G204gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n251_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT66), .A3(new_n259_), .ZN(new_n260_));
  OR3_X1    g059(.A1(new_n251_), .A2(KEYINPUT66), .A3(new_n257_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT13), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G229gat), .A2(G233gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT14), .ZN(new_n267_));
  AND2_X1   g066(.A1(KEYINPUT73), .A2(G1gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(KEYINPUT73), .A2(G1gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n267_), .B1(new_n270_), .B2(G8gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(G15gat), .B(G22gat), .Z(new_n272_));
  NOR3_X1   g071(.A1(new_n271_), .A2(KEYINPUT74), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT74), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT73), .B(G1gat), .ZN(new_n275_));
  INV_X1    g074(.A(G8gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT14), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n272_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n274_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(G1gat), .B1(new_n273_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT74), .B1(new_n271_), .B2(new_n272_), .ZN(new_n281_));
  INV_X1    g080(.A(G1gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n280_), .A2(G8gat), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(G8gat), .B1(new_n280_), .B2(new_n284_), .ZN(new_n286_));
  INV_X1    g085(.A(G29gat), .ZN(new_n287_));
  INV_X1    g086(.A(G36gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G43gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G29gat), .A2(G36gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G50gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n290_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G43gat), .ZN(new_n298_));
  AOI21_X1  g097(.A(G50gat), .B1(new_n298_), .B2(new_n292_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n285_), .A2(new_n286_), .A3(new_n301_), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n273_), .A2(new_n279_), .A3(G1gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n282_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n276_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n280_), .A2(G8gat), .A3(new_n284_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n300_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n266_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT15), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n294_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n298_), .A2(G50gat), .A3(new_n292_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(KEYINPUT15), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n305_), .A2(new_n300_), .A3(new_n306_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n265_), .A3(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G113gat), .B(G141gat), .ZN(new_n318_));
  INV_X1    g117(.A(G169gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G197gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n308_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT80), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n308_), .A2(KEYINPUT80), .A3(new_n317_), .A4(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n308_), .A2(new_n317_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n322_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n264_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G231gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n242_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(new_n306_), .A3(new_n305_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G183gat), .B(G211gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G155gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n343_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT17), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT77), .B1(new_n347_), .B2(KEYINPUT75), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT17), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n349_), .A3(new_n345_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(KEYINPUT77), .A3(new_n350_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n339_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n346_), .A2(KEYINPUT75), .A3(KEYINPUT17), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n337_), .A2(new_n355_), .A3(new_n338_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(KEYINPUT78), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT78), .B1(new_n354_), .B2(new_n356_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  OR2_X1    g162(.A1(G141gat), .A2(G148gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT86), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n364_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n368_), .B(KEYINPUT2), .Z(new_n369_));
  OAI211_X1 g168(.A(new_n362_), .B(new_n363_), .C1(new_n367_), .C2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n363_), .B(KEYINPUT1), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n368_), .B(new_n364_), .C1(new_n371_), .C2(new_n361_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  OR3_X1    g172(.A1(new_n373_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT28), .B1(new_n373_), .B2(KEYINPUT29), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G22gat), .B(G50gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n321_), .A2(G204gat), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n255_), .A2(G197gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT21), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n255_), .A3(G197gat), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT87), .B1(new_n321_), .B2(G204gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n385_), .B1(new_n386_), .B2(new_n380_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n382_), .B(new_n383_), .C1(new_n387_), .C2(KEYINPUT21), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT88), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n383_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n387_), .A2(new_n391_), .A3(KEYINPUT21), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n373_), .A2(KEYINPUT29), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G228gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n396_), .A3(new_n394_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(KEYINPUT89), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT89), .B1(new_n398_), .B2(new_n399_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n379_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G78gat), .B(G106gat), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n403_), .B(new_n405_), .C1(new_n401_), .C2(new_n379_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n379_), .A2(new_n401_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n402_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n378_), .B1(new_n408_), .B2(new_n400_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n404_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT83), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT31), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n414_), .B(new_n415_), .Z(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G127gat), .B(G134gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G113gat), .B(G120gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n419_), .B(new_n420_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(new_n418_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT30), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G176gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n319_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G169gat), .A2(G176gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(KEYINPUT24), .A3(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT81), .B(G190gat), .Z(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n431_), .B2(KEYINPUT26), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT25), .B(G183gat), .Z(new_n433_));
  OAI21_X1  g232(.A(new_n429_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n434_), .A2(KEYINPUT82), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G183gat), .A2(G190gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT23), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(KEYINPUT24), .B2(new_n427_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(KEYINPUT82), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n437_), .B1(G183gat), .B2(new_n431_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(G169gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n425_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n424_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n417_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT84), .B(G15gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n447_), .A2(new_n448_), .A3(new_n417_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n450_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n453_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n412_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n446_), .A2(new_n393_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n429_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n438_), .B2(KEYINPUT90), .ZN(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT26), .B(G190gat), .Z(new_n463_));
  OAI221_X1 g262(.A(new_n462_), .B1(KEYINPUT90), .B2(new_n438_), .C1(new_n433_), .C2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n437_), .B1(G183gat), .B2(G190gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT22), .B(G169gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT91), .Z(new_n467_));
  OAI211_X1 g266(.A(new_n428_), .B(new_n465_), .C1(new_n467_), .C2(G176gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n460_), .B(KEYINPUT20), .C1(new_n393_), .C2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G226gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT19), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n446_), .A2(new_n393_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n469_), .A2(new_n393_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n475_), .A2(KEYINPUT20), .A3(new_n472_), .A4(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT18), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(G64gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(new_n214_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT92), .B1(new_n478_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n482_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT92), .ZN(new_n485_));
  INV_X1    g284(.A(new_n482_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n474_), .A2(new_n485_), .A3(new_n477_), .A4(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT93), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G1gat), .B(G29gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(G85gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT0), .ZN(new_n492_));
  INV_X1    g291(.A(G57gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n373_), .A2(new_n423_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n370_), .A2(new_n422_), .A3(new_n372_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT96), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G225gat), .A2(G233gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(KEYINPUT4), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT94), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n501_), .B(new_n502_), .C1(KEYINPUT4), .C2(new_n495_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n502_), .B2(new_n501_), .ZN(new_n504_));
  AOI211_X1 g303(.A(new_n494_), .B(new_n500_), .C1(new_n504_), .C2(new_n499_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n499_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n497_), .A2(new_n499_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n494_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(KEYINPUT33), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n507_), .A2(new_n494_), .A3(new_n508_), .A4(new_n511_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n505_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT93), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n483_), .A2(new_n484_), .A3(new_n516_), .A4(new_n487_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n489_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  AND4_X1   g317(.A1(KEYINPUT20), .A2(new_n475_), .A3(new_n473_), .A4(new_n476_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(new_n472_), .B2(new_n470_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT97), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n482_), .A2(KEYINPUT32), .ZN(new_n522_));
  OR3_X1    g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n507_), .A2(new_n508_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n494_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n509_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n478_), .A2(new_n522_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n521_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n523_), .A2(new_n527_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n459_), .B1(new_n518_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n527_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n406_), .A2(new_n457_), .A3(new_n410_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n457_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT27), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n488_), .A2(new_n536_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n484_), .B(KEYINPUT27), .C1(new_n520_), .C2(new_n482_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n333_), .B(new_n360_), .C1(new_n531_), .C2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n314_), .A2(new_n234_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT69), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n234_), .A2(new_n301_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n314_), .A2(KEYINPUT69), .A3(new_n234_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT68), .B(KEYINPUT35), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .A4(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT67), .Z(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT34), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n544_), .A2(KEYINPUT70), .A3(new_n545_), .A4(new_n546_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n547_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT71), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G134gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(G162gat), .Z(new_n562_));
  AND2_X1   g361(.A1(new_n562_), .A2(KEYINPUT36), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(KEYINPUT36), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n554_), .B1(new_n552_), .B2(new_n556_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n558_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n552_), .A2(new_n556_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n553_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n564_), .B1(new_n569_), .B2(new_n557_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n541_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(G1gat), .B1(new_n574_), .B2(new_n532_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n575_), .A2(KEYINPUT98), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(KEYINPUT98), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n531_), .A2(new_n540_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n333_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT79), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n359_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(KEYINPUT79), .A3(new_n357_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT72), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT72), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n586_), .B(new_n587_), .C1(new_n567_), .C2(new_n570_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n569_), .B(new_n557_), .C1(new_n564_), .C2(new_n563_), .ZN(new_n589_));
  OAI22_X1  g388(.A1(new_n558_), .A2(new_n566_), .B1(KEYINPUT36), .B2(new_n562_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(KEYINPUT72), .A4(new_n585_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n584_), .A2(new_n588_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n578_), .A2(new_n579_), .A3(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n594_), .A2(new_n527_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT38), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n595_), .A2(new_n596_), .A3(new_n275_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n595_), .B2(new_n275_), .ZN(new_n598_));
  OAI22_X1  g397(.A1(new_n576_), .A2(new_n577_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT99), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT99), .ZN(new_n601_));
  OAI221_X1 g400(.A(new_n601_), .B1(new_n597_), .B2(new_n598_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(G1324gat));
  NAND3_X1  g402(.A1(new_n594_), .A2(new_n276_), .A3(new_n539_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n573_), .A2(new_n539_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n606_), .B2(G8gat), .ZN(new_n607_));
  AOI211_X1 g406(.A(KEYINPUT39), .B(new_n276_), .C1(new_n573_), .C2(new_n539_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g409(.A(G15gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n573_), .B2(new_n457_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT41), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n594_), .A2(new_n611_), .A3(new_n457_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1326gat));
  INV_X1    g414(.A(G22gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n594_), .A2(new_n616_), .A3(new_n411_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n573_), .A2(new_n411_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(G22gat), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n541_), .A2(new_n572_), .A3(new_n412_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT101), .B1(new_n621_), .B2(new_n616_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT100), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n620_), .A2(new_n625_), .A3(new_n622_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n624_), .A2(KEYINPUT42), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT42), .B1(new_n624_), .B2(new_n626_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n617_), .B1(new_n627_), .B2(new_n628_), .ZN(G1327gat));
  AND2_X1   g428(.A1(new_n518_), .A2(new_n530_), .ZN(new_n630_));
  OAI22_X1  g429(.A1(new_n630_), .A2(new_n459_), .B1(new_n539_), .B2(new_n535_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n584_), .A2(new_n571_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n631_), .A2(KEYINPUT102), .A3(new_n333_), .A4(new_n632_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n333_), .B(new_n632_), .C1(new_n531_), .C2(new_n540_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n287_), .A3(new_n527_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n588_), .A2(new_n591_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n531_), .B2(new_n540_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n584_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT43), .B(new_n639_), .C1(new_n531_), .C2(new_n540_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n642_), .A2(new_n333_), .A3(new_n643_), .A4(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT44), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n645_), .A2(new_n646_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n532_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n638_), .B1(new_n650_), .B2(new_n287_), .ZN(G1328gat));
  INV_X1    g450(.A(KEYINPUT46), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n645_), .B(KEYINPUT44), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n288_), .B1(new_n653_), .B2(new_n539_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n633_), .A2(new_n636_), .A3(new_n288_), .A4(new_n539_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT45), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n652_), .B1(new_n654_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n539_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n648_), .A2(new_n649_), .A3(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT46), .B(new_n656_), .C1(new_n660_), .C2(new_n288_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(G1329gat));
  NAND3_X1  g461(.A1(new_n633_), .A2(new_n636_), .A3(new_n457_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(KEYINPUT103), .A2(G43gat), .ZN(new_n664_));
  OR2_X1    g463(.A1(KEYINPUT103), .A2(G43gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n663_), .A2(KEYINPUT104), .A3(new_n664_), .A4(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n649_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n671_), .A2(G43gat), .A3(new_n457_), .A4(new_n647_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT47), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT47), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n670_), .A2(new_n672_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1330gat));
  NAND3_X1  g476(.A1(new_n637_), .A2(new_n294_), .A3(new_n411_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n648_), .A2(new_n649_), .A3(new_n412_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(new_n294_), .ZN(G1331gat));
  NOR2_X1   g479(.A1(new_n578_), .A2(new_n331_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n264_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n682_), .A2(new_n572_), .A3(new_n643_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n684_), .A2(new_n493_), .A3(new_n532_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n592_), .A2(new_n264_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT105), .Z(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(new_n681_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n688_), .A2(KEYINPUT106), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(KEYINPUT106), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n527_), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n691_), .B2(new_n493_), .ZN(G1332gat));
  INV_X1    g491(.A(G64gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n683_), .B2(new_n539_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n689_), .A2(new_n690_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n539_), .A2(new_n693_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n697_), .B2(new_n698_), .ZN(G1333gat));
  OAI21_X1  g498(.A(G71gat), .B1(new_n684_), .B2(new_n458_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(KEYINPUT49), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(KEYINPUT49), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n458_), .A2(G71gat), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT107), .Z(new_n704_));
  OAI22_X1  g503(.A1(new_n701_), .A2(new_n702_), .B1(new_n697_), .B2(new_n704_), .ZN(G1334gat));
  INV_X1    g504(.A(G78gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n683_), .B2(new_n411_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT50), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n411_), .A2(new_n706_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n697_), .B2(new_n710_), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n263_), .A2(new_n331_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .A4(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n713_), .A2(new_n213_), .A3(new_n532_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n682_), .A2(new_n571_), .A3(new_n584_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n527_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n716_), .B2(new_n213_), .ZN(G1336gat));
  NOR3_X1   g516(.A1(new_n713_), .A2(new_n214_), .A3(new_n659_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n539_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n214_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1337gat));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(KEYINPUT51), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n715_), .A2(new_n204_), .A3(new_n457_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G99gat), .B1(new_n713_), .B2(new_n458_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n723_), .A2(KEYINPUT51), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(G1338gat));
  OR2_X1    g528(.A1(new_n713_), .A2(new_n412_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n730_), .A2(G106gat), .A3(new_n731_), .A4(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n713_), .A2(new_n412_), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n732_), .B(new_n733_), .C1(new_n736_), .C2(new_n205_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n715_), .A2(new_n205_), .A3(new_n411_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n735_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT53), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT53), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n735_), .A2(new_n737_), .A3(new_n741_), .A4(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1339gat));
  INV_X1    g542(.A(G113gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT115), .B1(new_n332_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT57), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n246_), .A2(new_n203_), .A3(new_n248_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n246_), .A2(new_n248_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n202_), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT55), .B(new_n203_), .C1(new_n246_), .C2(new_n248_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(KEYINPUT56), .A3(new_n256_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  INV_X1    g555(.A(new_n747_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n749_), .A2(new_n202_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT55), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n249_), .A2(new_n748_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n756_), .B1(new_n761_), .B2(new_n257_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n752_), .A2(KEYINPUT111), .A3(KEYINPUT56), .A4(new_n256_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n755_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n258_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n265_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n315_), .A2(new_n266_), .A3(new_n316_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n767_), .A2(new_n322_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n764_), .A2(new_n766_), .B1(new_n262_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n746_), .B1(new_n771_), .B2(new_n572_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n764_), .A2(new_n766_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n262_), .A2(new_n770_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT57), .B(new_n571_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n762_), .A2(new_n778_), .A3(new_n753_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n752_), .B2(new_n256_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n765_), .B1(new_n780_), .B2(KEYINPUT113), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(new_n781_), .A3(new_n770_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n779_), .A2(new_n781_), .A3(new_n770_), .A4(KEYINPUT58), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n639_), .A3(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT112), .B(new_n746_), .C1(new_n771_), .C2(new_n572_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n774_), .A2(new_n777_), .A3(new_n786_), .A4(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n360_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n584_), .A2(new_n588_), .A3(new_n332_), .A4(new_n591_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT54), .B1(new_n264_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n592_), .A2(new_n792_), .A3(new_n332_), .A4(new_n263_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n788_), .A2(new_n789_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n539_), .A2(new_n532_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n533_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT59), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n777_), .A2(new_n786_), .A3(new_n772_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n799_), .A2(new_n643_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n800_));
  OR3_X1    g599(.A1(new_n800_), .A2(KEYINPUT59), .A3(new_n796_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n797_), .A2(new_n798_), .A3(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n798_), .B1(new_n797_), .B2(new_n801_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n745_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n794_), .A2(new_n332_), .A3(new_n796_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n745_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n803_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n797_), .A2(new_n798_), .A3(new_n801_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n806_), .A2(new_n744_), .B1(new_n810_), .B2(KEYINPUT115), .ZN(G1340gat));
  NAND3_X1  g610(.A1(new_n797_), .A2(new_n264_), .A3(new_n801_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G120gat), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n794_), .A2(new_n796_), .ZN(new_n814_));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n263_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n814_), .B(new_n816_), .C1(KEYINPUT60), .C2(new_n815_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n813_), .A2(new_n817_), .ZN(G1341gat));
  AOI21_X1  g617(.A(G127gat), .B1(new_n814_), .B2(new_n584_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n789_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g620(.A(G134gat), .B1(new_n814_), .B2(new_n572_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n639_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n824_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g624(.A1(new_n795_), .A2(new_n534_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT116), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n788_), .A2(new_n789_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n793_), .A2(new_n791_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT118), .B1(new_n832_), .B2(new_n332_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n794_), .A2(new_n827_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n331_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n833_), .A2(new_n834_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n835_), .B2(new_n331_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n794_), .A2(new_n827_), .A3(KEYINPUT118), .A4(new_n332_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT117), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G141gat), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n838_), .A2(new_n841_), .A3(G141gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1344gat));
  NAND2_X1  g645(.A1(new_n835_), .A2(new_n264_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT119), .B(G148gat), .Z(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1345gat));
  NAND2_X1  g648(.A1(new_n835_), .A2(new_n584_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT61), .B(G155gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1346gat));
  AOI21_X1  g651(.A(G162gat), .B1(new_n835_), .B2(new_n572_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n639_), .A2(G162gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT120), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n835_), .B2(new_n855_), .ZN(G1347gat));
  NOR2_X1   g655(.A1(new_n659_), .A2(new_n527_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n533_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n799_), .A2(new_n643_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n830_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n467_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n331_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT121), .B1(new_n860_), .B2(new_n331_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  NOR4_X1   g666(.A1(new_n800_), .A2(new_n867_), .A3(new_n332_), .A4(new_n858_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n865_), .B1(new_n869_), .B2(G169gat), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n866_), .A2(new_n868_), .A3(KEYINPUT62), .A4(new_n319_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n864_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT123), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n864_), .B(new_n874_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1348gat));
  XNOR2_X1  g675(.A(new_n860_), .B(KEYINPUT122), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n426_), .B1(new_n877_), .B2(new_n263_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n858_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n831_), .A2(G176gat), .A3(new_n264_), .A4(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1349gat));
  NAND3_X1  g682(.A1(new_n862_), .A2(new_n433_), .A3(new_n360_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n884_), .A2(KEYINPUT125), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(KEYINPUT125), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n794_), .A2(new_n858_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G183gat), .B1(new_n887_), .B2(new_n584_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n885_), .A2(new_n886_), .A3(new_n888_), .ZN(G1350gat));
  OAI21_X1  g688(.A(G190gat), .B1(new_n877_), .B2(new_n823_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n571_), .A2(new_n463_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n877_), .B2(new_n891_), .ZN(G1351gat));
  NOR3_X1   g691(.A1(new_n794_), .A2(new_n457_), .A3(new_n412_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n857_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n321_), .B1(new_n894_), .B2(new_n332_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n895_), .A2(KEYINPUT126), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n895_), .A2(KEYINPUT126), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n894_), .A2(new_n321_), .A3(new_n332_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(G1352gat));
  NOR2_X1   g698(.A1(new_n894_), .A2(new_n263_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n255_), .ZN(G1353gat));
  NOR2_X1   g700(.A1(new_n894_), .A2(new_n789_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n902_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT63), .B(G211gat), .Z(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n902_), .B2(new_n904_), .ZN(G1354gat));
  INV_X1    g704(.A(new_n894_), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n906_), .A2(G218gat), .A3(new_n639_), .ZN(new_n907_));
  AOI21_X1  g706(.A(G218gat), .B1(new_n906_), .B2(new_n572_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1355gat));
endmodule


