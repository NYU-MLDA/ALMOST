//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n956_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G127gat), .B(G134gat), .Z(new_n203_));
  XOR2_X1   g002(.A(G113gat), .B(G120gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT80), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT2), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n213_), .A2(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT81), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(KEYINPUT81), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT82), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n218_), .A2(new_n223_), .A3(KEYINPUT82), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n211_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n210_), .B(KEYINPUT1), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n209_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n217_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n212_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n206_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n211_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n218_), .A2(new_n223_), .A3(KEYINPUT82), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT82), .B1(new_n218_), .B2(new_n223_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n230_), .A2(new_n231_), .A3(new_n212_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n205_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(KEYINPUT4), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n238_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n206_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G1gat), .B(G29gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G57gat), .B(G85gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n246_), .B1(new_n233_), .B2(new_n239_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n247_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT96), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n245_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n252_), .B1(new_n258_), .B2(new_n254_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n247_), .A2(KEYINPUT96), .A3(new_n253_), .A4(new_n255_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT98), .Z(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT29), .B1(new_n228_), .B2(new_n232_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT85), .ZN(new_n265_));
  INV_X1    g064(.A(G197gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n266_), .B2(G204gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT84), .B(G197gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(G204gat), .ZN(new_n269_));
  INV_X1    g068(.A(G204gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT84), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(G197gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n266_), .A2(KEYINPUT84), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n265_), .B(new_n270_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n269_), .A2(KEYINPUT21), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT21), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n266_), .A2(KEYINPUT84), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(G197gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n270_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G197gat), .A2(G204gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n276_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G211gat), .B(G218gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n275_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT86), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n280_), .ZN(new_n286_));
  OAI211_X1 g085(.A(KEYINPUT86), .B(new_n286_), .C1(new_n268_), .C2(new_n270_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n282_), .A2(new_n276_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n283_), .A2(KEYINPUT87), .A3(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT87), .B1(new_n283_), .B2(new_n289_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n264_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G228gat), .A2(G233gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n269_), .A2(KEYINPUT21), .A3(new_n274_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n277_), .A2(new_n278_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n280_), .B1(new_n297_), .B2(G204gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n282_), .B1(new_n298_), .B2(KEYINPUT21), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n289_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n293_), .B(KEYINPUT83), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n264_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G78gat), .B(G106gat), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(KEYINPUT88), .Z(new_n306_));
  NAND3_X1  g105(.A1(new_n295_), .A2(new_n306_), .A3(new_n302_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G22gat), .B(G50gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT28), .B1(new_n241_), .B2(KEYINPUT29), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n241_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n310_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  OR3_X1    g113(.A1(new_n241_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(new_n311_), .A3(new_n309_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n305_), .A2(new_n308_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n306_), .B1(new_n295_), .B2(new_n302_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n317_), .B1(new_n308_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT89), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n317_), .B(KEYINPUT89), .C1(new_n308_), .C2(new_n319_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n318_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G169gat), .ZN(new_n325_));
  INV_X1    g124(.A(G176gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(KEYINPUT24), .ZN(new_n328_));
  INV_X1    g127(.A(G183gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT25), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT25), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G183gat), .ZN(new_n332_));
  INV_X1    g131(.A(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT26), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT26), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G190gat), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n330_), .A2(new_n332_), .A3(new_n334_), .A4(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n328_), .B1(new_n337_), .B2(KEYINPUT74), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT23), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(G183gat), .A3(G190gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n339_), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT25), .B(G183gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT26), .B(G190gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT24), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n351_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n327_), .A2(KEYINPUT75), .A3(KEYINPUT24), .A4(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n338_), .A2(new_n346_), .A3(new_n350_), .A4(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n325_), .A2(KEYINPUT22), .ZN(new_n359_));
  AOI21_X1  g158(.A(G176gat), .B1(new_n359_), .B2(KEYINPUT77), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT22), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(G169gat), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n363_), .B2(KEYINPUT77), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n340_), .A2(new_n342_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n329_), .A2(new_n333_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n341_), .A2(KEYINPUT78), .A3(G183gat), .A4(G190gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(new_n369_), .A3(new_n352_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n358_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G43gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n371_), .B(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(G15gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT30), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT79), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n374_), .A2(new_n379_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n384_));
  OR3_X1    g183(.A1(new_n383_), .A2(new_n384_), .A3(new_n205_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n205_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n324_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389_));
  XOR2_X1   g188(.A(G8gat), .B(G36gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT18), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n359_), .A2(new_n362_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT90), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n359_), .A2(new_n362_), .A3(KEYINPUT90), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n326_), .A3(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n344_), .A2(new_n367_), .A3(new_n345_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n352_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n328_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n327_), .A2(KEYINPUT24), .A3(new_n352_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n401_), .A2(new_n368_), .A3(new_n366_), .A4(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n300_), .A2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n283_), .A2(new_n358_), .A3(new_n289_), .A4(new_n370_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(KEYINPUT20), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT19), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT91), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n407_), .A2(KEYINPUT91), .A3(new_n409_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n409_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n371_), .B2(new_n300_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n418_));
  INV_X1    g217(.A(new_n300_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n404_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n300_), .A2(new_n404_), .A3(KEYINPUT92), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n415_), .B(new_n417_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n393_), .B1(new_n414_), .B2(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n407_), .A2(KEYINPUT91), .A3(new_n409_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT91), .B1(new_n407_), .B2(new_n409_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n393_), .B(new_n423_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n389_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n393_), .ZN(new_n430_));
  OR3_X1    g229(.A1(new_n290_), .A2(new_n291_), .A3(new_n404_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n415_), .B1(new_n431_), .B2(new_n417_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n407_), .A2(new_n409_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n430_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(new_n427_), .A3(KEYINPUT27), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n429_), .A2(new_n435_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n263_), .A2(new_n388_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n259_), .A2(KEYINPUT95), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n259_), .A2(KEYINPUT95), .A3(KEYINPUT33), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT93), .B1(new_n424_), .B2(new_n428_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n423_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n430_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT93), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n427_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n233_), .A2(new_n246_), .A3(new_n239_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n253_), .B(new_n448_), .C1(new_n244_), .C2(new_n246_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n442_), .A2(new_n443_), .A3(new_n447_), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n393_), .A2(KEYINPUT32), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n414_), .A2(new_n423_), .A3(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(KEYINPUT32), .B(new_n393_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT97), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n261_), .A4(new_n260_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n453_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT97), .B1(new_n262_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n324_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n324_), .A2(new_n436_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n262_), .B(KEYINPUT98), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n387_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n437_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G29gat), .B(G36gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G43gat), .B(G50gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT15), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT9), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G85gat), .B(G92gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT10), .B(G99gat), .ZN(new_n473_));
  OAI22_X1  g272(.A1(new_n471_), .A2(new_n472_), .B1(new_n473_), .B2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT64), .B(G85gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(G92gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n472_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n486_));
  INV_X1    g285(.A(G99gat), .ZN(new_n487_));
  INV_X1    g286(.A(G106gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n485_), .B1(new_n491_), .B2(new_n483_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n475_), .A2(new_n484_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT66), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n479_), .A2(KEYINPUT65), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n480_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n489_), .A2(KEYINPUT66), .A3(new_n490_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n499_), .A3(KEYINPUT6), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n496_), .A2(new_n501_), .A3(new_n502_), .A4(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n472_), .A2(new_n493_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n494_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n470_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G232gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT34), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT35), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n494_), .A2(new_n469_), .A3(new_n506_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n508_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n511_), .A2(new_n512_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G190gat), .B(G218gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G134gat), .B(G162gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(KEYINPUT36), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n515_), .A2(new_n516_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n515_), .A2(new_n516_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n520_), .B(KEYINPUT36), .Z(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n523_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G1gat), .B(G8gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT70), .B(G15gat), .Z(new_n533_));
  INV_X1    g332(.A(G22gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT70), .B(G15gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(G22gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(G8gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n532_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  AOI211_X1 g341(.A(new_n531_), .B(new_n542_), .C1(new_n535_), .C2(new_n537_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G71gat), .B(G78gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT11), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n548_));
  INV_X1    g347(.A(new_n546_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n547_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n544_), .B(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n553_), .A2(new_n555_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n557_), .A2(KEYINPUT17), .A3(new_n562_), .A4(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n562_), .B(KEYINPUT17), .Z(new_n565_));
  INV_X1    g364(.A(new_n563_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n565_), .B1(new_n566_), .B2(new_n556_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n552_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n505_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n502_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT66), .B1(new_n489_), .B2(new_n490_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n503_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT6), .B1(new_n497_), .B2(new_n499_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n570_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n489_), .A2(new_n490_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n481_), .A2(new_n482_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n472_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n579_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n581_));
  OAI22_X1  g380(.A1(new_n580_), .A2(KEYINPUT8), .B1(new_n581_), .B2(new_n474_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n569_), .B1(new_n577_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT12), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT12), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n507_), .A2(new_n585_), .A3(new_n569_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n494_), .A2(new_n506_), .A3(new_n552_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT67), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT67), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(new_n592_), .A3(new_n589_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n583_), .A2(new_n588_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n589_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT5), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G176gat), .B(G204gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n585_), .B1(new_n507_), .B2(new_n569_), .ZN(new_n605_));
  AOI211_X1 g404(.A(KEYINPUT12), .B(new_n552_), .C1(new_n494_), .C2(new_n506_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n593_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n592_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n597_), .B(new_n602_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n604_), .A2(KEYINPUT68), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT68), .ZN(new_n611_));
  INV_X1    g410(.A(new_n609_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n602_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n611_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n610_), .A2(new_n614_), .A3(KEYINPUT13), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT13), .B1(new_n610_), .B2(new_n614_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n469_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n537_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n536_), .A2(G22gat), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n540_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n531_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n538_), .A2(new_n532_), .A3(new_n540_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n469_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT73), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n621_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G229gat), .A2(G233gat), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT73), .B(new_n620_), .C1(new_n541_), .C2(new_n543_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n470_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n630_), .B(new_n627_), .C1(new_n634_), .C2(new_n544_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G113gat), .B(G141gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G169gat), .B(G197gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n637_), .B(new_n638_), .Z(new_n639_));
  XNOR2_X1  g438(.A(new_n636_), .B(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n619_), .A2(new_n641_), .ZN(new_n642_));
  NOR4_X1   g441(.A1(new_n466_), .A2(new_n530_), .A3(new_n568_), .A4(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n202_), .B1(new_n643_), .B2(new_n263_), .ZN(new_n644_));
  XOR2_X1   g443(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n645_));
  AND3_X1   g444(.A1(new_n517_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n527_), .B(KEYINPUT69), .Z(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n517_), .B2(new_n522_), .ZN(new_n648_));
  OAI21_X1  g447(.A(KEYINPUT37), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT37), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n523_), .B(new_n650_), .C1(new_n526_), .C2(new_n528_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n568_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT72), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n466_), .A2(new_n656_), .A3(new_n640_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n202_), .A3(new_n263_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n644_), .B1(new_n645_), .B2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n645_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n660_), .A2(KEYINPUT100), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(KEYINPUT100), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(G1324gat));
  NAND3_X1  g462(.A1(new_n657_), .A2(new_n539_), .A3(new_n436_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n643_), .A2(new_n436_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(G8gat), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT39), .B(new_n539_), .C1(new_n643_), .C2(new_n436_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n669_), .B(new_n670_), .Z(G1325gat));
  NAND3_X1  g470(.A1(new_n657_), .A2(new_n376_), .A3(new_n387_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n643_), .A2(new_n387_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n673_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(new_n673_), .B2(G15gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1326gat));
  INV_X1    g477(.A(new_n324_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n534_), .B1(new_n643_), .B2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n657_), .A2(new_n534_), .A3(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n466_), .A2(new_n640_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n653_), .A2(new_n529_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n619_), .A2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G29gat), .B1(new_n688_), .B2(new_n263_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n642_), .A2(new_n653_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n388_), .A2(new_n436_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n462_), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n459_), .A2(new_n324_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n387_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  INV_X1    g494(.A(new_n652_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT44), .B(new_n690_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n690_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n466_), .B2(new_n652_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT104), .B1(new_n704_), .B2(KEYINPUT44), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n690_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n700_), .B1(new_n705_), .B2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n263_), .A2(G29gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n689_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n685_), .A2(new_n713_), .A3(new_n436_), .A4(new_n687_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n699_), .A2(new_n436_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n705_), .B2(new_n709_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n718_), .B2(new_n713_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT46), .B(new_n716_), .C1(new_n718_), .C2(new_n713_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  NAND2_X1  g522(.A1(new_n387_), .A2(G43gat), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n724_), .B(new_n700_), .C1(new_n705_), .C2(new_n709_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n688_), .A2(new_n387_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT106), .B(G43gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT47), .B1(new_n725_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n724_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n710_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n728_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1330gat));
  AOI21_X1  g534(.A(G50gat), .B1(new_n688_), .B2(new_n679_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n679_), .A2(G50gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n710_), .B2(new_n737_), .ZN(G1331gat));
  NOR2_X1   g537(.A1(new_n466_), .A2(new_n530_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n619_), .A2(new_n641_), .A3(new_n568_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n462_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n619_), .A2(new_n641_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n694_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n568_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(G57gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n263_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n743_), .A2(new_n749_), .ZN(G1332gat));
  INV_X1    g549(.A(G64gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n741_), .B2(new_n436_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT48), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n747_), .A2(new_n751_), .A3(new_n436_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1333gat));
  INV_X1    g554(.A(G71gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n741_), .B2(new_n387_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT107), .B(KEYINPUT49), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n747_), .A2(new_n756_), .A3(new_n387_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1334gat));
  INV_X1    g560(.A(G78gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n741_), .B2(new_n679_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT50), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n747_), .A2(new_n762_), .A3(new_n679_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1335gat));
  NAND2_X1  g565(.A1(new_n702_), .A2(new_n703_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n702_), .A2(KEYINPUT108), .A3(new_n703_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n744_), .A2(new_n568_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n773_), .A2(new_n462_), .A3(new_n476_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n745_), .A2(new_n686_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G85gat), .B1(new_n775_), .B2(new_n263_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1336gat));
  INV_X1    g576(.A(new_n436_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G92gat), .B1(new_n773_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(G92gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n775_), .A2(new_n780_), .A3(new_n436_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1337gat));
  OAI21_X1  g581(.A(G99gat), .B1(new_n773_), .B2(new_n465_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n465_), .A2(new_n473_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n775_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT51), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n783_), .A2(new_n788_), .A3(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1338gat));
  NAND3_X1  g589(.A1(new_n775_), .A2(new_n488_), .A3(new_n679_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n771_), .A2(new_n324_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n767_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n794_), .B2(G106gat), .ZN(new_n795_));
  AOI211_X1 g594(.A(KEYINPUT52), .B(new_n488_), .C1(new_n767_), .C2(new_n793_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n791_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n797_), .B(new_n799_), .ZN(G1339gat));
  NOR2_X1   g599(.A1(new_n640_), .A2(new_n612_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n587_), .A2(KEYINPUT55), .A3(new_n591_), .A4(new_n593_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n588_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n596_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n803_), .A2(new_n804_), .A3(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n807_), .A2(KEYINPUT56), .A3(new_n603_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT56), .B1(new_n807_), .B2(new_n603_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n801_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n639_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n636_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n634_), .A2(new_n544_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n627_), .A2(new_n631_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n629_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n811_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n817_), .B2(KEYINPUT112), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(new_n819_), .A3(new_n811_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n812_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n610_), .A2(new_n614_), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n530_), .B1(new_n810_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT57), .B1(new_n823_), .B2(KEYINPUT113), .ZN(new_n824_));
  INV_X1    g623(.A(new_n636_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n639_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n609_), .B1(new_n826_), .B2(new_n812_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n807_), .A2(new_n603_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n807_), .A2(KEYINPUT56), .A3(new_n603_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n827_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n610_), .A2(new_n614_), .A3(new_n821_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n529_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n824_), .A2(new_n837_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n594_), .A2(new_n802_), .B1(new_n596_), .B2(new_n805_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n602_), .B1(new_n839_), .B2(new_n804_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT116), .B1(new_n840_), .B2(KEYINPUT56), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n831_), .A2(KEYINPUT115), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n828_), .A2(new_n843_), .A3(new_n829_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n807_), .A2(new_n845_), .A3(KEYINPUT56), .A4(new_n603_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n841_), .A2(new_n842_), .A3(new_n844_), .A4(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n818_), .A2(new_n820_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n812_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n609_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n821_), .A2(KEYINPUT114), .A3(new_n609_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT58), .B1(new_n847_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n847_), .A2(new_n854_), .A3(KEYINPUT58), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n696_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n653_), .B1(new_n838_), .B2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n746_), .B(new_n640_), .C1(new_n615_), .C2(new_n617_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT54), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT111), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n655_), .A2(KEYINPUT110), .A3(new_n864_), .A4(new_n640_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n860_), .A2(KEYINPUT111), .A3(KEYINPUT54), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT110), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n860_), .B2(KEYINPUT54), .ZN(new_n868_));
  AND4_X1   g667(.A1(new_n863_), .A2(new_n865_), .A3(new_n866_), .A4(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n263_), .B(new_n691_), .C1(new_n859_), .C2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(G113gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n641_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n870_), .A2(new_n875_), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n847_), .A2(KEYINPUT58), .A3(new_n854_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n877_), .A2(new_n855_), .A3(new_n652_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n824_), .A2(new_n837_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n568_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n863_), .A2(new_n865_), .A3(new_n866_), .A4(new_n868_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n462_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT59), .B1(new_n882_), .B2(new_n691_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n874_), .B1(new_n876_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n870_), .A2(new_n875_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n882_), .A2(KEYINPUT59), .A3(new_n691_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(KEYINPUT117), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n640_), .B1(new_n884_), .B2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n873_), .B1(new_n888_), .B2(new_n872_), .ZN(G1340gat));
  AOI21_X1  g688(.A(new_n619_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n890_));
  INV_X1    g689(.A(G120gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n619_), .B2(KEYINPUT60), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(KEYINPUT60), .B2(new_n891_), .ZN(new_n893_));
  OAI22_X1  g692(.A1(new_n890_), .A2(new_n891_), .B1(new_n870_), .B2(new_n893_), .ZN(G1341gat));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT119), .B(G127gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n653_), .A2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n884_), .B2(new_n887_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n880_), .A2(new_n881_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n899_), .A2(new_n263_), .A3(new_n691_), .A4(new_n653_), .ZN(new_n900_));
  INV_X1    g699(.A(G127gat), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT118), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n900_), .A2(new_n904_), .A3(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n895_), .B1(new_n898_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n897_), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n885_), .A2(KEYINPUT117), .A3(new_n886_), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT117), .B1(new_n885_), .B2(new_n886_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n903_), .A2(new_n905_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n912_), .A3(KEYINPUT120), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n907_), .A2(new_n913_), .ZN(G1342gat));
  INV_X1    g713(.A(G134gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n871_), .A2(new_n915_), .A3(new_n530_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n652_), .B1(new_n884_), .B2(new_n887_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n915_), .ZN(G1343gat));
  NOR3_X1   g717(.A1(new_n324_), .A2(new_n387_), .A3(new_n436_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n882_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n641_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g722(.A(new_n619_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n921_), .A2(new_n924_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g725(.A1(new_n920_), .A2(new_n568_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT61), .B(G155gat), .Z(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1346gat));
  INV_X1    g728(.A(G162gat), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n920_), .A2(new_n930_), .A3(new_n652_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n920_), .B2(new_n529_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n933_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n931_), .B1(new_n934_), .B2(new_n935_), .ZN(G1347gat));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n462_), .A2(new_n436_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n388_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n899_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n640_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n937_), .B1(new_n942_), .B2(G169gat), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n396_), .A2(new_n397_), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n943_), .A2(new_n944_), .B1(new_n945_), .B2(new_n941_), .ZN(new_n946_));
  OR2_X1    g745(.A1(new_n943_), .A2(new_n944_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n941_), .A2(KEYINPUT122), .A3(new_n325_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n946_), .B1(new_n947_), .B2(new_n948_), .ZN(G1348gat));
  INV_X1    g748(.A(new_n940_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n950_), .B(new_n924_), .C1(new_n951_), .C2(G176gat), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(G176gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(KEYINPUT124), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n952_), .B(new_n954_), .ZN(G1349gat));
  NOR2_X1   g754(.A1(new_n940_), .A2(new_n568_), .ZN(new_n956_));
  MUX2_X1   g755(.A(G183gat), .B(new_n347_), .S(new_n956_), .Z(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n940_), .B2(new_n652_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n530_), .A2(new_n348_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n940_), .B2(new_n959_), .ZN(G1351gat));
  NOR3_X1   g759(.A1(new_n938_), .A2(new_n324_), .A3(new_n387_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n899_), .A2(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n962_), .A2(new_n640_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(new_n266_), .ZN(G1352gat));
  NAND3_X1  g763(.A1(new_n899_), .A2(new_n924_), .A3(new_n961_), .ZN(new_n965_));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  NAND4_X1  g766(.A1(new_n899_), .A2(KEYINPUT125), .A3(new_n924_), .A4(new_n961_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n967_), .A2(G204gat), .A3(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n970_));
  INV_X1    g769(.A(new_n965_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n970_), .B1(new_n971_), .B2(new_n270_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n969_), .A2(new_n972_), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974_));
  NAND4_X1  g773(.A1(new_n967_), .A2(new_n970_), .A3(G204gat), .A4(new_n968_), .ZN(new_n975_));
  AND3_X1   g774(.A1(new_n973_), .A2(new_n974_), .A3(new_n975_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n974_), .B1(new_n973_), .B2(new_n975_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n976_), .A2(new_n977_), .ZN(G1353gat));
  NOR2_X1   g777(.A1(new_n962_), .A2(new_n568_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n980_));
  AND2_X1   g779(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n979_), .B1(new_n980_), .B2(new_n981_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n982_), .B1(new_n979_), .B2(new_n980_), .ZN(G1354gat));
  OAI21_X1  g782(.A(G218gat), .B1(new_n962_), .B2(new_n652_), .ZN(new_n984_));
  OR2_X1    g783(.A1(new_n529_), .A2(G218gat), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n984_), .B1(new_n962_), .B2(new_n985_), .ZN(G1355gat));
endmodule


