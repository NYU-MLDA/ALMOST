//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  XOR2_X1   g004(.A(G127gat), .B(G134gat), .Z(new_n206_));
  XOR2_X1   g005(.A(G113gat), .B(G120gat), .Z(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT83), .Z(new_n210_));
  INV_X1    g009(.A(G155gat), .ZN(new_n211_));
  INV_X1    g010(.A(G162gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G141gat), .ZN(new_n215_));
  INV_X1    g014(.A(G148gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT2), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n217_), .A2(new_n219_), .B1(new_n221_), .B2(KEYINPUT3), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT84), .B(KEYINPUT3), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n223_), .A2(KEYINPUT85), .A3(new_n221_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT85), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT84), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT84), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT3), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n225_), .B1(new_n230_), .B2(new_n220_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n222_), .B1(new_n224_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT85), .B1(new_n223_), .B2(new_n221_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n225_), .A3(new_n220_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(KEYINPUT86), .A3(new_n222_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n214_), .B1(new_n234_), .B2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n215_), .A2(new_n216_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n209_), .B(KEYINPUT83), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n241_), .A2(KEYINPUT1), .B1(new_n211_), .B2(new_n212_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n210_), .A2(new_n243_), .ZN(new_n244_));
  AOI211_X1 g043(.A(new_n220_), .B(new_n240_), .C1(new_n242_), .C2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n208_), .B1(new_n239_), .B2(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n237_), .A2(KEYINPUT86), .A3(new_n222_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT86), .B1(new_n237_), .B2(new_n222_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n213_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n242_), .A2(new_n244_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n240_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n221_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n208_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G225gat), .A2(G233gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n246_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n246_), .A2(KEYINPUT4), .A3(new_n254_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n258_), .B(new_n208_), .C1(new_n239_), .C2(new_n245_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n255_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n205_), .B(new_n256_), .C1(new_n257_), .C2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT96), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(KEYINPUT33), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n246_), .A2(KEYINPUT4), .A3(new_n254_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(new_n260_), .A3(new_n259_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n268_), .A2(new_n205_), .A3(new_n256_), .A4(new_n264_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n259_), .A2(new_n255_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT97), .B1(new_n257_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT97), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n267_), .A2(new_n272_), .A3(new_n255_), .A4(new_n259_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n246_), .A2(new_n254_), .A3(new_n260_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n205_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n266_), .A2(new_n269_), .B1(new_n274_), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT18), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G64gat), .B(G92gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(G169gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT22), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT22), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G169gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT93), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n285_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n283_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(KEYINPUT80), .A2(G183gat), .A3(G190gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT23), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n293_), .A2(KEYINPUT23), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n292_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n300_), .B(KEYINPUT92), .Z(new_n301_));
  NAND3_X1  g100(.A1(new_n291_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT26), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(G190gat), .ZN(new_n304_));
  INV_X1    g103(.A(G190gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(KEYINPUT26), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT91), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT25), .B(G183gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(KEYINPUT26), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n303_), .A2(G190gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT91), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n307_), .A2(new_n308_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(new_n284_), .A3(new_n283_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n315_), .A2(KEYINPUT24), .A3(new_n316_), .A4(new_n300_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n316_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT24), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n295_), .A2(new_n296_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(new_n322_), .B2(KEYINPUT23), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n313_), .A2(new_n317_), .A3(new_n320_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n302_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G197gat), .B(G204gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT21), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(G197gat), .A2(G204gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G197gat), .A2(G204gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(KEYINPUT21), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G211gat), .B(G218gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n331_), .A2(new_n332_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n325_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n323_), .A2(new_n292_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(G169gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n317_), .B(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n320_), .B(new_n344_), .C1(new_n298_), .C2(new_n297_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n335_), .B(new_n341_), .C1(new_n343_), .C2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n337_), .A2(KEYINPUT20), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n348_), .A3(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n341_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n336_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n335_), .A2(new_n302_), .A3(new_n324_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n355_), .A2(KEYINPUT20), .A3(new_n351_), .A4(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n348_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n282_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT95), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n347_), .A2(new_n352_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT94), .ZN(new_n363_));
  INV_X1    g162(.A(new_n282_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(new_n357_), .A4(new_n353_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(KEYINPUT95), .B(new_n282_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n268_), .A2(new_n256_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n276_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n262_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n354_), .A2(new_n336_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n356_), .A2(KEYINPUT20), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n352_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n337_), .A2(new_n346_), .A3(KEYINPUT20), .A4(new_n351_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT98), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n363_), .A2(new_n357_), .A3(new_n353_), .A4(new_n377_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n376_), .A2(KEYINPUT98), .A3(new_n378_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n278_), .A2(new_n368_), .B1(new_n371_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n249_), .A2(new_n386_), .A3(new_n252_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT28), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT28), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n249_), .A2(new_n389_), .A3(new_n386_), .A4(new_n252_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G22gat), .B(G50gat), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT89), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G228gat), .ZN(new_n395_));
  INV_X1    g194(.A(G233gat), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n396_), .A2(KEYINPUT87), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(KEYINPUT87), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT88), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G78gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n399_), .B(KEYINPUT88), .ZN(new_n403_));
  INV_X1    g202(.A(G78gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G106gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n234_), .A2(new_n238_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n245_), .B1(new_n408_), .B2(new_n213_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n336_), .B1(new_n409_), .B2(new_n386_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n407_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n391_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n389_), .B1(new_n409_), .B2(new_n386_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n390_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n394_), .A2(new_n411_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n416_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n407_), .A2(new_n410_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n407_), .A2(new_n410_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n419_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT99), .B1(new_n385_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n266_), .A2(new_n269_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n274_), .A2(new_n277_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n368_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n384_), .A2(new_n371_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT99), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n419_), .A2(new_n423_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n371_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n366_), .A2(new_n367_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n376_), .B2(new_n282_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n365_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n425_), .A2(new_n433_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT100), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(G43gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n354_), .B(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(G15gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT30), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n445_), .B(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT81), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n208_), .B(KEYINPUT31), .Z(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n449_), .A2(KEYINPUT81), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n453_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT82), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(KEYINPUT82), .A3(new_n455_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n441_), .A2(new_n442_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n442_), .B1(new_n441_), .B2(new_n460_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT101), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n439_), .A2(new_n463_), .A3(new_n432_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n436_), .A2(new_n438_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT101), .B1(new_n465_), .B2(new_n424_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n456_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(new_n371_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n461_), .A2(new_n462_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G229gat), .A2(G233gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G1gat), .B(G8gat), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G1gat), .A2(G8gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT14), .ZN(new_n476_));
  AND2_X1   g275(.A1(G15gat), .A2(G22gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(G15gat), .A2(G22gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT71), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n479_), .A2(KEYINPUT71), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT72), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n482_), .A2(KEYINPUT72), .A3(new_n483_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n474_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n473_), .A3(new_n484_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n472_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n487_), .A2(new_n489_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n492_), .B(KEYINPUT15), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n493_), .A3(new_n471_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G113gat), .B(G141gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT76), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G169gat), .B(G197gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT77), .B1(new_n501_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT77), .ZN(new_n507_));
  INV_X1    g306(.A(new_n505_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n496_), .A2(new_n500_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n501_), .A2(new_n505_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n470_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G231gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(new_n396_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n497_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n497_), .A2(new_n517_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n524_));
  XOR2_X1   g323(.A(G71gat), .B(G78gat), .Z(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT67), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT67), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n521_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n519_), .A2(new_n520_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G127gat), .B(G155gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G183gat), .B(G211gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n542_), .A2(KEYINPUT17), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(KEYINPUT17), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n537_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT74), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n537_), .A2(KEYINPUT74), .A3(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n521_), .A2(new_n528_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n528_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n534_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n543_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT34), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT35), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(G85gat), .ZN(new_n563_));
  INV_X1    g362(.A(G92gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568_));
  NOR2_X1   g367(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT6), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n567_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT66), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT66), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n576_), .B(new_n567_), .C1(new_n570_), .C2(new_n573_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n575_), .A2(KEYINPUT8), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT8), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(KEYINPUT66), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n565_), .A2(new_n581_), .A3(new_n566_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n565_), .A2(new_n566_), .B1(new_n581_), .B2(G92gat), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT64), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n583_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT64), .B1(new_n582_), .B2(new_n584_), .ZN(new_n588_));
  INV_X1    g387(.A(G106gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT10), .B(G99gat), .Z(new_n590_));
  AOI21_X1  g389(.A(new_n573_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n587_), .A2(new_n588_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n580_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n578_), .A2(new_n593_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n594_), .A2(new_n492_), .B1(new_n559_), .B2(new_n558_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT68), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n578_), .B2(new_n593_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n575_), .A2(KEYINPUT8), .A3(new_n577_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n598_), .A2(KEYINPUT68), .A3(new_n580_), .A4(new_n592_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n599_), .A3(new_n498_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n562_), .B1(new_n595_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n560_), .A2(new_n561_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n603_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n603_), .A2(new_n608_), .ZN(new_n611_));
  OR3_X1    g410(.A1(new_n610_), .A2(new_n611_), .A3(KEYINPUT37), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT37), .B1(new_n610_), .B2(new_n611_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n555_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n535_), .B1(new_n578_), .B2(new_n593_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n594_), .A2(new_n532_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n552_), .A2(KEYINPUT12), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n597_), .A2(new_n599_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT69), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n597_), .A2(new_n599_), .A3(KEYINPUT69), .A4(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n617_), .A2(KEYINPUT12), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n623_), .A2(new_n624_), .B1(new_n625_), .B2(new_n616_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n618_), .B1(new_n626_), .B2(new_n615_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT5), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n629_), .B(new_n630_), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n627_), .B(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(KEYINPUT13), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(KEYINPUT13), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n614_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT75), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n514_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n371_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n639_), .A2(G1gat), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n424_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n440_), .B1(new_n648_), .B2(new_n431_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n385_), .A2(KEYINPUT99), .A3(new_n424_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n460_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT100), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n441_), .A2(new_n442_), .A3(new_n460_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n469_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n610_), .A2(new_n611_), .A3(KEYINPUT103), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT103), .B1(new_n610_), .B2(new_n611_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n555_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n635_), .A2(new_n513_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n640_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n643_), .A2(new_n644_), .A3(KEYINPUT38), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n647_), .A2(new_n665_), .A3(new_n666_), .ZN(G1324gat));
  OR3_X1    g466(.A1(new_n639_), .A2(G8gat), .A3(new_n439_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n663_), .A2(new_n465_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(G8gat), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(G8gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT40), .Z(G1325gat));
  NOR3_X1   g473(.A1(new_n639_), .A2(G15gat), .A3(new_n460_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT105), .ZN(new_n676_));
  OAI21_X1  g475(.A(G15gat), .B1(new_n664_), .B2(new_n460_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT41), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(KEYINPUT41), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n676_), .A2(new_n678_), .A3(new_n679_), .ZN(G1326gat));
  INV_X1    g479(.A(G22gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n663_), .B2(new_n424_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n424_), .A2(new_n681_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n639_), .B2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(new_n658_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n555_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n687_), .A2(new_n635_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n514_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n371_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n662_), .A2(new_n688_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n612_), .A2(new_n613_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n469_), .B1(new_n651_), .B2(KEYINPUT100), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT43), .B(new_n694_), .C1(new_n695_), .C2(new_n653_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  INV_X1    g496(.A(new_n694_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n655_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n693_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n470_), .B2(new_n694_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n655_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(KEYINPUT44), .A3(new_n693_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n702_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n371_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n692_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  NAND3_X1  g508(.A1(new_n702_), .A2(new_n706_), .A3(new_n465_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n439_), .A2(G36gat), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n655_), .A2(new_n512_), .A3(new_n689_), .A4(new_n712_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n713_), .A2(KEYINPUT107), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(KEYINPUT107), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(KEYINPUT45), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT45), .B1(new_n714_), .B2(new_n715_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n711_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n711_), .A2(KEYINPUT46), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  NAND4_X1  g522(.A1(new_n702_), .A2(new_n706_), .A3(G43gat), .A4(new_n467_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n690_), .A2(new_n460_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(G43gat), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n691_), .B2(new_n424_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n424_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n707_), .B2(new_n729_), .ZN(G1331gat));
  NAND2_X1  g529(.A1(new_n614_), .A2(new_n635_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT108), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n732_), .A2(new_n512_), .A3(new_n470_), .ZN(new_n733_));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n371_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n635_), .A2(new_n513_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT109), .B1(new_n660_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n738_));
  INV_X1    g537(.A(new_n736_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n655_), .A2(new_n738_), .A3(new_n659_), .A4(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n737_), .A2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(new_n371_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n735_), .B1(new_n742_), .B2(new_n734_), .ZN(G1332gat));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n733_), .A2(new_n744_), .A3(new_n465_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n741_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G64gat), .B1(new_n746_), .B2(new_n439_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(KEYINPUT48), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(KEYINPUT48), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1333gat));
  INV_X1    g549(.A(G71gat), .ZN(new_n751_));
  INV_X1    g550(.A(new_n460_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n733_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n737_), .A2(new_n752_), .A3(new_n740_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(G71gat), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G71gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(G1334gat));
  NAND3_X1  g559(.A1(new_n733_), .A2(new_n404_), .A3(new_n424_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G78gat), .B1(new_n746_), .B2(new_n432_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(KEYINPUT50), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(KEYINPUT50), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n736_), .A2(new_n688_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769_), .B2(new_n640_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n470_), .A2(new_n512_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n687_), .A2(new_n636_), .A3(new_n688_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n563_), .A3(new_n371_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n775_), .ZN(G1336gat));
  OAI21_X1  g575(.A(G92gat), .B1(new_n769_), .B2(new_n439_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n564_), .A3(new_n465_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1337gat));
  NAND2_X1  g578(.A1(new_n768_), .A2(new_n752_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G99gat), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n467_), .A2(new_n590_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n773_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT113), .ZN(new_n786_));
  NAND2_X1  g585(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n781_), .A2(new_n789_), .A3(new_n784_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n792_));
  AOI211_X1 g591(.A(KEYINPUT113), .B(new_n783_), .C1(new_n780_), .C2(G99gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n787_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(G1338gat));
  AOI211_X1 g594(.A(new_n432_), .B(new_n767_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n589_), .B1(new_n796_), .B2(KEYINPUT115), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n424_), .B(new_n766_), .C1(new_n696_), .C2(new_n699_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT52), .B1(new_n797_), .B2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n705_), .A2(KEYINPUT115), .A3(new_n424_), .A4(new_n766_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n800_), .A2(new_n802_), .A3(KEYINPUT52), .A4(G106gat), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n771_), .A2(new_n589_), .A3(new_n424_), .A4(new_n772_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT114), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n801_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n802_), .A2(G106gat), .ZN(new_n809_));
  INV_X1    g608(.A(new_n800_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n803_), .A4(new_n805_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n807_), .A2(new_n813_), .ZN(G1339gat));
  NAND3_X1  g613(.A1(new_n614_), .A2(new_n636_), .A3(new_n513_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n623_), .A2(new_n624_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n625_), .A2(new_n616_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n615_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n824_), .A3(new_n822_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n626_), .A2(KEYINPUT55), .A3(new_n615_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT116), .B1(new_n626_), .B2(new_n615_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n823_), .A2(new_n825_), .A3(new_n826_), .A4(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n631_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n828_), .A2(KEYINPUT56), .A3(new_n631_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(KEYINPUT119), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n631_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n825_), .A2(new_n827_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n626_), .A2(KEYINPUT55), .A3(new_n615_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT55), .B1(new_n626_), .B2(new_n615_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n834_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(KEYINPUT56), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n471_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n499_), .A2(new_n493_), .A3(new_n472_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n505_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT118), .B1(new_n510_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n510_), .A2(KEYINPUT118), .A3(new_n844_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n846_), .A2(new_n847_), .B1(new_n627_), .B2(new_n834_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n833_), .A2(new_n841_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n694_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n848_), .A4(new_n841_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n627_), .A2(new_n834_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n847_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n845_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT56), .B1(new_n828_), .B2(new_n631_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n840_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n859_), .B2(new_n832_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n860_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n841_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n851_), .A2(new_n854_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n632_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n839_), .B2(KEYINPUT56), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n858_), .A2(KEYINPUT117), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n832_), .A3(new_n867_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n512_), .A2(new_n855_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n864_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n863_), .B1(new_n870_), .B2(new_n658_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n832_), .B1(new_n858_), .B2(KEYINPUT117), .ZN(new_n872_));
  AOI211_X1 g671(.A(new_n865_), .B(KEYINPUT56), .C1(new_n828_), .C2(new_n631_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n869_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n864_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(KEYINPUT57), .A3(new_n687_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n862_), .A2(new_n871_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n817_), .B1(new_n878_), .B2(new_n555_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n468_), .A2(new_n640_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n882_), .A2(KEYINPUT59), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(KEYINPUT59), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n513_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(G113gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT121), .B1(new_n879_), .B2(new_n881_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n876_), .B2(new_n687_), .ZN(new_n889_));
  AOI211_X1 g688(.A(new_n863_), .B(new_n658_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n688_), .B1(new_n891_), .B2(new_n862_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n888_), .B(new_n880_), .C1(new_n892_), .C2(new_n817_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n887_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n512_), .A2(new_n886_), .ZN(new_n895_));
  OAI22_X1  g694(.A1(new_n885_), .A2(new_n886_), .B1(new_n894_), .B2(new_n895_), .ZN(G1340gat));
  AOI21_X1  g695(.A(new_n636_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n897_));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n636_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(KEYINPUT60), .B2(new_n898_), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n897_), .A2(new_n898_), .B1(new_n894_), .B2(new_n900_), .ZN(G1341gat));
  AOI21_X1  g700(.A(new_n555_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n902_));
  INV_X1    g701(.A(G127gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n688_), .A2(new_n903_), .ZN(new_n904_));
  OAI22_X1  g703(.A1(new_n902_), .A2(new_n903_), .B1(new_n894_), .B2(new_n904_), .ZN(G1342gat));
  INV_X1    g704(.A(G134gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n694_), .A2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT123), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n887_), .A2(new_n893_), .A3(new_n658_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n906_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n910_), .A2(KEYINPUT122), .A3(new_n906_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n909_), .B1(new_n913_), .B2(new_n914_), .ZN(G1343gat));
  NOR4_X1   g714(.A1(new_n752_), .A2(new_n432_), .A3(new_n640_), .A4(new_n465_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n892_), .B2(new_n817_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n513_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n215_), .ZN(G1344gat));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n636_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n216_), .ZN(G1345gat));
  NOR2_X1   g720(.A1(new_n917_), .A2(new_n555_), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT61), .B(G155gat), .Z(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1346gat));
  OAI21_X1  g723(.A(G162gat), .B1(new_n917_), .B2(new_n694_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n658_), .A2(new_n212_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n917_), .B2(new_n926_), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n879_), .A2(new_n439_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n460_), .A2(new_n424_), .A3(new_n371_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n928_), .A2(new_n512_), .A3(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n930_), .A2(new_n931_), .A3(G169gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n928_), .A2(new_n929_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n934_), .B(new_n512_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n931_), .B1(new_n930_), .B2(G169gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n932_), .B1(new_n935_), .B2(new_n936_), .ZN(G1348gat));
  NOR2_X1   g736(.A1(new_n933_), .A2(new_n636_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n283_), .ZN(G1349gat));
  AOI21_X1  g738(.A(G183gat), .B1(new_n934_), .B2(new_n688_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n933_), .A2(new_n308_), .A3(new_n555_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n933_), .B2(new_n694_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n658_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n933_), .B2(new_n944_), .ZN(G1351gat));
  AND2_X1   g744(.A1(new_n460_), .A2(new_n434_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n928_), .A2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n512_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n636_), .B1(new_n950_), .B2(G204gat), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n947_), .A2(new_n951_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n950_), .A2(G204gat), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n952_), .B(new_n954_), .ZN(G1353gat));
  NOR3_X1   g754(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956_));
  AOI211_X1 g755(.A(new_n956_), .B(new_n555_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n947_), .A2(new_n957_), .ZN(new_n958_));
  OAI21_X1  g757(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(KEYINPUT126), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n958_), .B(new_n960_), .ZN(G1354gat));
  NAND2_X1  g760(.A1(new_n947_), .A2(new_n658_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(KEYINPUT127), .B(G218gat), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n694_), .A2(new_n963_), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n962_), .A2(new_n963_), .B1(new_n947_), .B2(new_n964_), .ZN(G1355gat));
endmodule


