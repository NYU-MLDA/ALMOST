//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n917_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202_));
  XOR2_X1   g001(.A(G1gat), .B(G29gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT99), .B(G85gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT0), .B(G57gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT98), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT4), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT80), .ZN(new_n211_));
  INV_X1    g010(.A(G127gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(G134gat), .ZN(new_n213_));
  INV_X1    g012(.A(G134gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(G127gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n211_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(G127gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(G134gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT80), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G113gat), .B(G120gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n220_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT80), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT80), .B1(new_n217_), .B2(new_n218_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G141gat), .ZN(new_n226_));
  INV_X1    g025(.A(G148gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT81), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G155gat), .A3(G162gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n232_), .B1(new_n237_), .B2(KEYINPUT1), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n234_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n231_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n229_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n232_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n221_), .B(new_n225_), .C1(new_n241_), .C2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT95), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n235_), .B1(G155gat), .B2(G162gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n233_), .A2(KEYINPUT81), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT1), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n232_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n240_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n230_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n225_), .A2(new_n221_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n248_), .A2(new_n249_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n251_), .A2(new_n252_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n260_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n259_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(KEYINPUT95), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n210_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT96), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G225gat), .A2(G233gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT97), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n251_), .B2(KEYINPUT4), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n263_), .A2(KEYINPUT97), .A3(new_n210_), .A4(new_n264_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n268_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n209_), .B1(new_n267_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n262_), .A2(new_n265_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT96), .B1(new_n274_), .B2(KEYINPUT4), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT96), .ZN(new_n276_));
  AOI211_X1 g075(.A(new_n276_), .B(new_n210_), .C1(new_n262_), .C2(new_n265_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n209_), .B(new_n272_), .C1(new_n275_), .C2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n268_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n208_), .B1(new_n273_), .B2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G197gat), .A2(G204gat), .ZN(new_n282_));
  INV_X1    g081(.A(G197gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT85), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G197gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n282_), .B1(new_n287_), .B2(G204gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT87), .B1(new_n288_), .B2(KEYINPUT21), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n290_), .B1(new_n283_), .B2(G204gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT85), .B(G197gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(G204gat), .ZN(new_n293_));
  INV_X1    g092(.A(G204gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n287_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n295_), .A3(KEYINPUT21), .ZN(new_n296_));
  INV_X1    g095(.A(new_n282_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT21), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n289_), .A2(new_n296_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n288_), .A2(KEYINPUT88), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT88), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n302_), .A2(new_n300_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n257_), .A2(new_n230_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT83), .B(G228gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT84), .B(G233gat), .ZN(new_n313_));
  OAI221_X1 g112(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT89), .B1(new_n311_), .B2(new_n310_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT89), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n316_), .B(KEYINPUT29), .C1(new_n241_), .C2(new_n250_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n309_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT90), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n312_), .A2(new_n313_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n319_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n314_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G78gat), .B(G106gat), .Z(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n324_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n314_), .B(new_n326_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n311_), .B2(new_n310_), .ZN(new_n330_));
  NOR4_X1   g129(.A1(new_n241_), .A2(new_n250_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT82), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n258_), .A2(new_n310_), .A3(new_n260_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT28), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n311_), .A2(new_n329_), .A3(new_n310_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G22gat), .B(G50gat), .Z(new_n338_));
  AND3_X1   g137(.A1(new_n332_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT91), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n332_), .A2(new_n337_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n338_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT91), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n332_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n328_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n347_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n272_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT98), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n353_), .A2(new_n207_), .A3(new_n279_), .A4(new_n278_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n281_), .A2(new_n349_), .A3(new_n351_), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT19), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n303_), .A2(new_n308_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT23), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(G183gat), .B2(G190gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT22), .B(G169gat), .Z(new_n362_));
  INV_X1    g161(.A(KEYINPUT92), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G169gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT92), .ZN(new_n366_));
  INV_X1    g165(.A(G176gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n368_), .A2(KEYINPUT93), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT93), .B1(new_n368_), .B2(new_n369_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n361_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n373_), .A2(G169gat), .A3(G176gat), .ZN(new_n374_));
  INV_X1    g173(.A(G169gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT77), .B1(new_n375_), .B2(new_n367_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n377_), .A2(KEYINPUT24), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT26), .B(G190gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT25), .B(G183gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(KEYINPUT24), .A3(new_n369_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n378_), .A2(new_n360_), .A3(new_n381_), .A4(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n358_), .B1(new_n372_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G183gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT25), .B1(new_n385_), .B2(KEYINPUT75), .ZN(new_n386_));
  OR3_X1    g185(.A1(new_n385_), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT26), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n389_), .A2(G190gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(G190gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n388_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n386_), .B(new_n387_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n394_), .A2(new_n378_), .A3(new_n360_), .A4(new_n382_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n369_), .B1(new_n362_), .B2(G176gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT78), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n398_), .B(new_n369_), .C1(new_n362_), .C2(G176gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n390_), .A2(new_n385_), .A3(new_n391_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n360_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n395_), .A2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT20), .B1(new_n309_), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n357_), .B1(new_n384_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n358_), .A2(new_n372_), .A3(new_n383_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT94), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n309_), .A2(new_n403_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n309_), .B2(new_n403_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n406_), .B(KEYINPUT20), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n405_), .B1(new_n410_), .B2(new_n357_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G8gat), .B(G36gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT18), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G64gat), .B(G92gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n405_), .B(new_n415_), .C1(new_n410_), .C2(new_n357_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT27), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n418_), .A2(KEYINPUT27), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n410_), .A2(new_n357_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n384_), .A2(new_n357_), .A3(new_n404_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n416_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n202_), .B1(new_n355_), .B2(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n281_), .A2(new_n354_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n349_), .A2(new_n351_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n420_), .A2(new_n419_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT103), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n354_), .A2(KEYINPUT33), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n278_), .A2(new_n279_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n207_), .A4(new_n353_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n268_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n267_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n207_), .B1(new_n274_), .B2(new_n438_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT100), .Z(new_n442_));
  AOI21_X1  g241(.A(new_n419_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n424_), .B1(new_n357_), .B2(new_n410_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n415_), .A2(KEYINPUT32), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT102), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT102), .ZN(new_n447_));
  INV_X1    g246(.A(new_n445_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n447_), .B(new_n448_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n445_), .B(KEYINPUT101), .Z(new_n450_));
  OR2_X1    g249(.A1(new_n411_), .A2(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n446_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n281_), .A2(new_n354_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n437_), .A2(new_n443_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n428_), .B(new_n432_), .C1(new_n454_), .C2(new_n430_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G227gat), .A2(G233gat), .ZN(new_n456_));
  INV_X1    g255(.A(G71gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(G99gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n403_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(new_n264_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G15gat), .B(G43gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT79), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT30), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT31), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n461_), .B(new_n465_), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n349_), .A2(new_n351_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n429_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n431_), .A2(new_n466_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT104), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n427_), .A2(new_n467_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT104), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n468_), .A4(new_n429_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n455_), .A2(new_n467_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G29gat), .B(G36gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G43gat), .B(G50gat), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT73), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485_));
  INV_X1    g284(.A(G1gat), .ZN(new_n486_));
  INV_X1    g285(.A(G8gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G1gat), .B(G8gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT74), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n484_), .A2(new_n491_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n482_), .B(KEYINPUT15), .ZN(new_n499_));
  INV_X1    g298(.A(new_n491_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n492_), .A2(new_n501_), .A3(new_n496_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G113gat), .B(G141gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(G169gat), .B(G197gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n503_), .B(new_n506_), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n475_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G120gat), .B(G148gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT5), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G176gat), .B(G204gat), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n511_), .B(new_n512_), .Z(new_n513_));
  XNOR2_X1  g312(.A(G85gat), .B(G92gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  INV_X1    g315(.A(G106gat), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n515_), .A2(KEYINPUT9), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT6), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G85gat), .A2(G92gat), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n518_), .B(new_n521_), .C1(KEYINPUT9), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT65), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(G99gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n517_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT64), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT7), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(new_n517_), .A3(KEYINPUT64), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n528_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n531_), .B1(G99gat), .B2(G106gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n535_), .A3(new_n527_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(new_n525_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT67), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(KEYINPUT65), .A3(new_n533_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT65), .B1(new_n530_), .B2(KEYINPUT7), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n536_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT67), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n539_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n538_), .A2(new_n543_), .A3(new_n521_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n524_), .B1(new_n544_), .B2(new_n515_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n515_), .A2(new_n524_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n521_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT66), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n539_), .A2(new_n541_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(KEYINPUT66), .A3(new_n521_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n546_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n523_), .B1(new_n545_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT11), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(KEYINPUT11), .ZN(new_n556_));
  XOR2_X1   g355(.A(G71gat), .B(G78gat), .Z(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n556_), .A2(new_n557_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n553_), .A2(new_n561_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n560_), .B(new_n523_), .C1(new_n545_), .C2(new_n552_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT68), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT68), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(new_n569_), .A3(new_n566_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n562_), .A2(KEYINPUT12), .A3(new_n563_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT12), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n553_), .A2(new_n573_), .A3(new_n561_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n566_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n513_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n574_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n565_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n513_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n578_), .A2(new_n568_), .A3(new_n570_), .A4(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT13), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n491_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(new_n560_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT16), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n587_), .A2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT72), .Z(new_n595_));
  AND2_X1   g394(.A1(new_n591_), .A2(new_n592_), .ZN(new_n596_));
  OR3_X1    g395(.A1(new_n587_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT37), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT34), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT35), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT70), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n553_), .B2(new_n499_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n603_), .A2(new_n604_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n520_), .B1(new_n550_), .B2(KEYINPUT67), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n514_), .B1(new_n611_), .B2(new_n543_), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n548_), .B(new_n520_), .C1(new_n541_), .C2(new_n539_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT66), .B1(new_n550_), .B2(new_n521_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI22_X1  g414(.A1(new_n524_), .A2(new_n612_), .B1(new_n615_), .B2(new_n546_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n616_), .A2(KEYINPUT69), .A3(new_n482_), .A4(new_n523_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n553_), .A2(new_n499_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT69), .ZN(new_n619_));
  INV_X1    g418(.A(new_n482_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n619_), .B1(new_n553_), .B2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n610_), .A2(new_n617_), .A3(new_n618_), .A4(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT71), .ZN(new_n624_));
  XOR2_X1   g423(.A(G134gat), .B(G162gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n621_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n499_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n616_), .B2(new_n523_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n608_), .B1(new_n631_), .B2(new_n606_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n628_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n627_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n622_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n622_), .B2(new_n633_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n600_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n622_), .A2(new_n633_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n634_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n622_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(KEYINPUT37), .A3(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n637_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n509_), .A2(new_n584_), .A3(new_n599_), .A4(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT105), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n486_), .A3(new_n453_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n640_), .A2(new_n641_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT106), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n475_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n584_), .A2(new_n507_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n598_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n654_), .B2(new_n429_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n646_), .A2(new_n647_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n648_), .A2(new_n655_), .A3(new_n656_), .ZN(G1324gat));
  NAND3_X1  g456(.A1(new_n645_), .A2(new_n487_), .A3(new_n427_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G8gat), .B1(new_n654_), .B2(new_n431_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT39), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(KEYINPUT39), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n658_), .B(KEYINPUT40), .C1(new_n660_), .C2(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1325gat));
  OAI21_X1  g465(.A(G15gat), .B1(new_n654_), .B2(new_n467_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT41), .Z(new_n668_));
  OR2_X1    g467(.A1(new_n467_), .A2(G15gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n644_), .B2(new_n669_), .ZN(G1326gat));
  OAI21_X1  g469(.A(G22gat), .B1(new_n654_), .B2(new_n468_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT42), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n468_), .A2(G22gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n644_), .B2(new_n673_), .ZN(G1327gat));
  OAI21_X1  g473(.A(KEYINPUT43), .B1(new_n475_), .B2(new_n643_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n432_), .A2(new_n428_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n437_), .A2(new_n443_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n452_), .A2(new_n453_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n430_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n467_), .B1(new_n676_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n471_), .A2(new_n474_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n637_), .A2(new_n642_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n675_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n584_), .A2(new_n507_), .A3(new_n598_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT44), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n690_), .B(new_n687_), .C1(new_n675_), .C2(new_n685_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n689_), .A2(new_n691_), .A3(new_n429_), .ZN(new_n692_));
  INV_X1    g491(.A(G29gat), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n649_), .B(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(new_n599_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n583_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n509_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n453_), .A2(new_n693_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT107), .ZN(new_n702_));
  OAI22_X1  g501(.A1(new_n692_), .A2(new_n693_), .B1(new_n700_), .B2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(G36gat), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n431_), .B(KEYINPUT109), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n699_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT45), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n689_), .A2(new_n691_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT108), .B1(new_n708_), .B2(new_n427_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n683_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT43), .B(new_n643_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n688_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n690_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n686_), .A2(KEYINPUT44), .A3(new_n688_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n713_), .A2(KEYINPUT108), .A3(new_n427_), .A4(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G36gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n707_), .B1(new_n709_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(KEYINPUT46), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  OAI221_X1 g519(.A(new_n707_), .B1(new_n718_), .B2(KEYINPUT46), .C1(new_n709_), .C2(new_n716_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  INV_X1    g521(.A(G43gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n699_), .A2(new_n723_), .A3(new_n466_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n689_), .A2(new_n691_), .A3(new_n467_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n723_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n699_), .B2(new_n430_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n430_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n708_), .B2(new_n730_), .ZN(G1331gat));
  NOR2_X1   g530(.A1(new_n475_), .A2(new_n507_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n643_), .A2(new_n599_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n584_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G57gat), .B1(new_n736_), .B2(new_n453_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n584_), .A2(new_n507_), .A3(new_n598_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n651_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(G57gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n453_), .B2(KEYINPUT111), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(KEYINPUT111), .B2(new_n741_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n737_), .B1(new_n740_), .B2(new_n743_), .ZN(G1332gat));
  INV_X1    g543(.A(G64gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n740_), .B2(new_n705_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT48), .Z(new_n747_));
  NAND2_X1  g546(.A1(new_n705_), .A2(new_n745_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT112), .Z(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n735_), .B2(new_n749_), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n739_), .B2(new_n467_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT49), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n736_), .A2(new_n457_), .A3(new_n466_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1334gat));
  OAI21_X1  g553(.A(G78gat), .B1(new_n739_), .B2(new_n468_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT50), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n468_), .A2(G78gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n735_), .B2(new_n757_), .ZN(G1335gat));
  NOR3_X1   g557(.A1(new_n584_), .A2(new_n507_), .A3(new_n599_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n686_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n429_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n732_), .A2(new_n583_), .A3(new_n696_), .ZN(new_n762_));
  OR3_X1    g561(.A1(new_n762_), .A2(G85gat), .A3(new_n429_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1336gat));
  INV_X1    g563(.A(new_n762_), .ZN(new_n765_));
  INV_X1    g564(.A(G92gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n427_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n686_), .A2(new_n705_), .A3(new_n759_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n766_), .ZN(G1337gat));
  NOR2_X1   g568(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n770_));
  OAI21_X1  g569(.A(G99gat), .B1(new_n760_), .B2(new_n467_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n765_), .A2(new_n466_), .A3(new_n516_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n773_), .B(new_n774_), .Z(G1338gat));
  NAND3_X1  g574(.A1(new_n765_), .A2(new_n517_), .A3(new_n430_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n686_), .A2(new_n430_), .A3(new_n759_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(G106gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n777_), .B2(G106gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g581(.A1(new_n470_), .A2(new_n430_), .A3(new_n429_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n572_), .A2(new_n566_), .A3(new_n574_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n786_), .A2(new_n575_), .A3(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n577_), .A2(new_n787_), .A3(new_n565_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n513_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n785_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n572_), .A2(new_n566_), .A3(new_n574_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n578_), .A2(KEYINPUT55), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n579_), .B1(new_n575_), .B2(new_n787_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT115), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(KEYINPUT56), .A3(new_n796_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT116), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n795_), .A2(new_n796_), .A3(new_n801_), .A4(KEYINPUT56), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n793_), .A2(new_n798_), .A3(new_n800_), .A4(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n507_), .A2(new_n580_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n498_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n495_), .A2(new_n496_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n496_), .B1(new_n484_), .B2(new_n491_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n506_), .B1(new_n808_), .B2(new_n501_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n806_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n581_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n581_), .A2(KEYINPUT117), .A3(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n805_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT57), .B1(new_n817_), .B2(new_n695_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n791_), .A2(new_n799_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n811_), .A2(new_n580_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n791_), .B2(new_n799_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT58), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n684_), .A3(new_n824_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n803_), .A2(new_n804_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n695_), .A2(KEYINPUT57), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n598_), .B1(new_n818_), .B2(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n733_), .A2(new_n583_), .A3(new_n507_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NOR4_X1   g634(.A1(new_n733_), .A2(new_n583_), .A3(new_n507_), .A4(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n784_), .B1(new_n829_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(G113gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n507_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n684_), .B1(new_n823_), .B2(KEYINPUT58), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n819_), .B(new_n821_), .C1(new_n791_), .C2(new_n799_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n650_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n817_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n845_), .B1(new_n826_), .B2(new_n650_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n599_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n830_), .A2(new_n834_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n841_), .B(new_n783_), .C1(new_n849_), .C2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n829_), .A2(new_n837_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n855_), .A2(KEYINPUT118), .A3(new_n841_), .A4(new_n783_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n783_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT59), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n857_), .A2(new_n507_), .A3(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n840_), .B1(new_n860_), .B2(new_n839_), .ZN(G1340gat));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n584_), .B1(new_n858_), .B2(KEYINPUT59), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n857_), .B2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n584_), .A2(KEYINPUT60), .ZN(new_n865_));
  MUX2_X1   g664(.A(KEYINPUT60), .B(new_n865_), .S(new_n862_), .Z(new_n866_));
  NAND2_X1  g665(.A1(new_n838_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT119), .B1(new_n864_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n583_), .B1(new_n838_), .B2(new_n841_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n870_), .B(new_n867_), .C1(new_n872_), .C2(new_n862_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n869_), .A2(new_n873_), .ZN(G1341gat));
  NAND3_X1  g673(.A1(new_n838_), .A2(new_n212_), .A3(new_n599_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n857_), .A2(new_n599_), .A3(new_n859_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n212_), .ZN(G1342gat));
  NAND3_X1  g676(.A1(new_n838_), .A2(new_n214_), .A3(new_n650_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n857_), .A2(new_n684_), .A3(new_n859_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n214_), .ZN(G1343gat));
  NOR4_X1   g679(.A1(new_n705_), .A2(new_n466_), .A3(new_n468_), .A4(new_n429_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT120), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n855_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n508_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT121), .B(G141gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1344gat));
  NOR2_X1   g685(.A1(new_n883_), .A2(new_n584_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n227_), .ZN(G1345gat));
  OR3_X1    g687(.A1(new_n883_), .A2(KEYINPUT122), .A3(new_n598_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT122), .B1(new_n883_), .B2(new_n598_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1346gat));
  INV_X1    g693(.A(new_n883_), .ZN(new_n895_));
  AOI21_X1  g694(.A(G162gat), .B1(new_n895_), .B2(new_n650_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n684_), .A2(G162gat), .ZN(new_n897_));
  XOR2_X1   g696(.A(new_n897_), .B(KEYINPUT123), .Z(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n895_), .B2(new_n898_), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n469_), .A2(new_n467_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n705_), .B(new_n900_), .C1(new_n849_), .C2(new_n851_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n901_), .A2(new_n508_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n364_), .A2(new_n366_), .ZN(new_n903_));
  OAI21_X1  g702(.A(G169gat), .B1(new_n901_), .B2(new_n508_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  OAI22_X1  g704(.A1(new_n902_), .A2(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n905_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT124), .B1(new_n906_), .B2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n902_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  OR3_X1    g710(.A1(new_n901_), .A2(new_n903_), .A3(new_n508_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n907_), .A4(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n909_), .A2(new_n913_), .ZN(G1348gat));
  NOR2_X1   g713(.A1(new_n901_), .A2(new_n584_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(new_n367_), .ZN(G1349gat));
  NOR2_X1   g715(.A1(new_n901_), .A2(new_n598_), .ZN(new_n917_));
  MUX2_X1   g716(.A(G183gat), .B(new_n380_), .S(new_n917_), .Z(G1350gat));
  NAND2_X1  g717(.A1(new_n650_), .A2(new_n379_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n901_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n921_), .B(G190gat), .C1(new_n901_), .C2(new_n643_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n855_), .A2(new_n684_), .A3(new_n705_), .A4(new_n900_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n921_), .B1(new_n924_), .B2(G190gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n920_), .B1(new_n923_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT126), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n928_), .B(new_n920_), .C1(new_n923_), .C2(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1351gat));
  NOR2_X1   g729(.A1(new_n355_), .A2(new_n466_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n855_), .A2(new_n705_), .A3(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n508_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n283_), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n584_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n294_), .ZN(G1353gat));
  NOR2_X1   g735(.A1(new_n932_), .A2(new_n598_), .ZN(new_n937_));
  OR2_X1    g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  XOR2_X1   g738(.A(KEYINPUT63), .B(G211gat), .Z(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(new_n937_), .B2(new_n940_), .ZN(G1354gat));
  OR3_X1    g740(.A1(new_n932_), .A2(G218gat), .A3(new_n695_), .ZN(new_n942_));
  OAI21_X1  g741(.A(G218gat), .B1(new_n932_), .B2(new_n643_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(KEYINPUT127), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n942_), .A2(new_n946_), .A3(new_n943_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1355gat));
endmodule


