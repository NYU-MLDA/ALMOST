//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G197gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(G197gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT21), .B1(new_n204_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT84), .B1(new_n203_), .B2(G204gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT84), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(new_n205_), .A3(G197gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n209_), .B(new_n211_), .C1(G197gat), .C2(new_n205_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n207_), .B(new_n208_), .C1(new_n212_), .C2(KEYINPUT21), .ZN(new_n213_));
  INV_X1    g012(.A(new_n208_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(KEYINPUT21), .A3(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT85), .ZN(new_n217_));
  AND2_X1   g016(.A1(G228gat), .A2(G233gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT80), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT80), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G141gat), .A3(G148gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n231_));
  NOR4_X1   g030(.A1(new_n231_), .A2(KEYINPUT81), .A3(G141gat), .A4(G148gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT3), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n229_), .B(new_n230_), .C1(new_n232_), .C2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT82), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n231_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(new_n234_), .A3(KEYINPUT3), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n223_), .B1(new_n237_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n222_), .B1(new_n221_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(new_n245_), .B2(new_n221_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n225_), .A2(new_n227_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n233_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n244_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT29), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n219_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G78gat), .ZN(new_n255_));
  INV_X1    g054(.A(G78gat), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n219_), .B(new_n256_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n218_), .A2(new_n217_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G22gat), .B(G50gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n252_), .A2(new_n253_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n262_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n265_), .A3(new_n261_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n258_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT86), .B(G106gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n268_), .A2(new_n258_), .A3(new_n270_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n273_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n274_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n276_), .B1(new_n277_), .B2(new_n271_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280_));
  INV_X1    g079(.A(G183gat), .ZN(new_n281_));
  INV_X1    g080(.A(G190gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285_));
  INV_X1    g084(.A(G169gat), .ZN(new_n286_));
  INV_X1    g085(.A(G176gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n283_), .A2(new_n284_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n287_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(KEYINPUT24), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G190gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n293_), .A2(KEYINPUT78), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT25), .B(G183gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT78), .B1(new_n282_), .B2(KEYINPUT26), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n289_), .B(new_n292_), .C1(new_n294_), .C2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n281_), .A2(new_n282_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n283_), .A2(new_n284_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G169gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT79), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n287_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n286_), .A2(KEYINPUT22), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n303_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n300_), .B(new_n291_), .C1(new_n305_), .C2(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n298_), .A2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT20), .B1(new_n309_), .B2(new_n216_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT19), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n300_), .A2(KEYINPUT89), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT89), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n283_), .A2(new_n315_), .A3(new_n284_), .A4(new_n299_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n291_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT22), .B(G169gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(new_n287_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n314_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT90), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT90), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n314_), .A2(new_n322_), .A3(new_n316_), .A4(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n291_), .A2(KEYINPUT24), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n324_), .A2(KEYINPUT88), .B1(new_n286_), .B2(new_n287_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(KEYINPUT88), .B2(new_n324_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n293_), .A2(new_n295_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n289_), .A2(new_n327_), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n321_), .A2(new_n323_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n216_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n313_), .A2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n298_), .A2(new_n213_), .A3(new_n215_), .A4(new_n308_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT20), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT87), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n321_), .A2(new_n323_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n328_), .A2(new_n326_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n216_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n335_), .A2(new_n336_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n312_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n331_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G8gat), .B(G36gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n332_), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT87), .B1(new_n332_), .B2(KEYINPUT20), .ZN(new_n351_));
  OAI22_X1  g150(.A1(new_n350_), .A2(new_n351_), .B1(new_n216_), .B2(new_n329_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n352_), .A2(new_n312_), .B1(new_n330_), .B2(new_n313_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n348_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n349_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n216_), .A2(new_n338_), .A3(new_n320_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n312_), .B1(new_n358_), .B2(new_n310_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n352_), .B2(new_n312_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n348_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n357_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n356_), .A2(new_n357_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G71gat), .B(G99gat), .ZN(new_n364_));
  INV_X1    g163(.A(G43gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n309_), .B(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G127gat), .B(G134gat), .Z(new_n368_));
  XOR2_X1   g167(.A(G113gat), .B(G120gat), .Z(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n367_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(G15gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT30), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT31), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n371_), .B(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n380_), .B(new_n370_), .C1(new_n244_), .C2(new_n251_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n237_), .A2(new_n243_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n223_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n370_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(new_n250_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n370_), .B1(new_n244_), .B2(new_n251_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n379_), .B(new_n381_), .C1(new_n388_), .C2(new_n380_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n378_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G1gat), .B(G29gat), .Z(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G57gat), .B(G85gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n386_), .A2(KEYINPUT4), .A3(new_n387_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n381_), .A2(new_n379_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n390_), .B(new_n396_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n377_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n279_), .A2(new_n363_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT96), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n279_), .A2(KEYINPUT96), .A3(new_n363_), .A4(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n402_), .ZN(new_n409_));
  AND4_X1   g208(.A1(new_n409_), .A2(new_n363_), .A3(new_n275_), .A4(new_n278_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n352_), .A2(new_n312_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n411_), .A2(new_n354_), .A3(new_n331_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n354_), .B1(new_n411_), .B2(new_n331_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n401_), .A2(KEYINPUT33), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT33), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n389_), .A2(new_n416_), .A3(new_n390_), .A4(new_n396_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n378_), .B(new_n381_), .C1(new_n388_), .C2(new_n380_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n378_), .B1(new_n388_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n386_), .A2(KEYINPUT93), .A3(new_n387_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n396_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n419_), .B1(new_n423_), .B2(KEYINPUT94), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n425_));
  AOI211_X1 g224(.A(new_n425_), .B(new_n396_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n414_), .B(new_n418_), .C1(new_n424_), .C2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT95), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n388_), .A2(new_n420_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n379_), .A3(new_n422_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n397_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n425_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n423_), .A2(KEYINPUT94), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n419_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n435_), .A2(KEYINPUT95), .A3(new_n414_), .A4(new_n418_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n343_), .B1(KEYINPUT32), .B2(new_n354_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n360_), .A2(KEYINPUT32), .A3(new_n354_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n402_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n429_), .A2(new_n436_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n410_), .B1(new_n441_), .B2(new_n279_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n377_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n408_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G99gat), .ZN(new_n448_));
  INV_X1    g247(.A(G106gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(KEYINPUT64), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT7), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT7), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n452_), .A2(new_n448_), .A3(new_n449_), .A4(KEYINPUT64), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n447_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G85gat), .ZN(new_n455_));
  INV_X1    g254(.A(G92gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G85gat), .A2(G92gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT65), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G36gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(G29gat), .ZN(new_n468_));
  INV_X1    g267(.A(G29gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(G36gat), .ZN(new_n470_));
  INV_X1    g269(.A(G50gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G43gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n365_), .A2(G50gat), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n468_), .A2(new_n470_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n468_), .A2(new_n470_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n454_), .A2(new_n464_), .A3(new_n460_), .ZN(new_n479_));
  OR2_X1    g278(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n449_), .A3(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n457_), .A2(KEYINPUT9), .A3(new_n458_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n458_), .A2(KEYINPUT9), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n447_), .A2(new_n482_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n466_), .A2(new_n478_), .A3(new_n479_), .A4(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G232gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT34), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n466_), .A2(new_n479_), .A3(new_n485_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT69), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT15), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n468_), .A2(new_n470_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n472_), .A2(new_n473_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(KEYINPUT15), .A3(new_n474_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n494_), .A2(new_n495_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n495_), .B1(new_n494_), .B2(new_n503_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n493_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n489_), .A2(new_n490_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G190gat), .B(G218gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT70), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G134gat), .B(G162gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n454_), .A2(new_n464_), .A3(new_n460_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n464_), .B1(new_n454_), .B2(new_n460_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n485_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT69), .B1(new_n518_), .B2(new_n502_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n494_), .A2(new_n495_), .A3(new_n503_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n507_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n493_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n508_), .A2(new_n514_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n508_), .A2(new_n523_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n512_), .B(new_n513_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n525_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  AOI211_X1 g328(.A(KEYINPUT72), .B(new_n527_), .C1(new_n508_), .C2(new_n523_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n524_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n444_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(G57gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(G64gat), .ZN(new_n534_));
  INV_X1    g333(.A(G64gat), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(G57gat), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT66), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(G57gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n533_), .A2(G64gat), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT66), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT11), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n537_), .A2(new_n544_), .A3(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n256_), .A2(G71gat), .ZN(new_n546_));
  INV_X1    g345(.A(G71gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(G78gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(new_n545_), .A3(new_n549_), .ZN(new_n550_));
  AOI211_X1 g349(.A(new_n544_), .B(new_n549_), .C1(new_n537_), .C2(new_n541_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(G8gat), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT73), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI211_X1 g356(.A(KEYINPUT73), .B(KEYINPUT14), .C1(new_n202_), .C2(new_n554_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G1gat), .B(G8gat), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n560_), .A2(new_n561_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n553_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT75), .ZN(new_n568_));
  XOR2_X1   g367(.A(G127gat), .B(G155gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(G183gat), .B(G211gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n568_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n567_), .A2(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT17), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n578_), .B1(new_n579_), .B2(new_n575_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n549_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n542_), .B2(KEYINPUT11), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n551_), .B1(new_n583_), .B2(new_n545_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n494_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n518_), .A2(new_n553_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n494_), .A2(new_n584_), .A3(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .A4(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n585_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n588_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT5), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G176gat), .B(G204gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n592_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT68), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n592_), .A2(KEYINPUT68), .A3(new_n595_), .A4(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n599_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT13), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT13), .ZN(new_n608_));
  AOI211_X1 g407(.A(new_n608_), .B(new_n605_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n564_), .A2(new_n478_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n477_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(KEYINPUT76), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT76), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n560_), .A2(new_n561_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n560_), .A2(new_n561_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n478_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n562_), .A2(new_n563_), .A3(new_n477_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n613_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n503_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n611_), .A3(new_n620_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT77), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G169gat), .B(G197gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n622_), .A2(new_n624_), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n610_), .A2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n532_), .A2(new_n581_), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n202_), .B1(new_n633_), .B2(new_n402_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT97), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n629_), .A2(new_n630_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n279_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n427_), .A2(new_n428_), .B1(new_n402_), .B2(new_n439_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(new_n436_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n377_), .B1(new_n639_), .B2(new_n410_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n636_), .B1(new_n640_), .B2(new_n408_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT37), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n642_), .B(new_n524_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT71), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n522_), .B1(new_n521_), .B2(new_n493_), .ZN(new_n645_));
  AOI211_X1 g444(.A(new_n507_), .B(new_n492_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n528_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n524_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n644_), .B1(new_n648_), .B2(KEYINPUT37), .ZN(new_n649_));
  AOI211_X1 g448(.A(KEYINPUT71), .B(new_n642_), .C1(new_n647_), .C2(new_n524_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n643_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n581_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n641_), .A2(new_n610_), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(new_n202_), .A3(new_n402_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT38), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n635_), .A2(new_n656_), .ZN(G1324gat));
  INV_X1    g456(.A(new_n363_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n554_), .B1(new_n633_), .B2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT39), .Z(new_n660_));
  NAND3_X1  g459(.A1(new_n654_), .A2(new_n554_), .A3(new_n658_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g462(.A(new_n373_), .B1(new_n633_), .B2(new_n443_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT41), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n654_), .A2(new_n373_), .A3(new_n443_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1326gat));
  INV_X1    g466(.A(G22gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n633_), .B2(new_n637_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT42), .Z(new_n670_));
  NAND3_X1  g469(.A1(new_n654_), .A2(new_n668_), .A3(new_n637_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n580_), .A2(new_n531_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n641_), .A2(new_n610_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n402_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n444_), .A2(new_n652_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT98), .B1(new_n676_), .B2(KEYINPUT43), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(KEYINPUT43), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT98), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n444_), .A2(new_n679_), .A3(new_n680_), .A4(new_n652_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n677_), .A2(new_n678_), .A3(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n632_), .A2(new_n580_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n683_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n684_), .A2(G29gat), .A3(new_n402_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT44), .B1(new_n682_), .B2(new_n683_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n675_), .B1(new_n685_), .B2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(KEYINPUT46), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n674_), .A2(new_n467_), .A3(new_n658_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT99), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n674_), .A2(new_n693_), .A3(new_n467_), .A4(new_n658_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT45), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n692_), .A2(new_n697_), .A3(new_n694_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n690_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n689_), .A2(KEYINPUT46), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n684_), .A2(new_n658_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G36gat), .B1(new_n701_), .B2(new_n686_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n699_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n700_), .B1(new_n699_), .B2(new_n702_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1329gat));
  NOR2_X1   g504(.A1(new_n377_), .A2(new_n365_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n684_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT101), .B1(new_n707_), .B2(new_n686_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n687_), .A2(new_n709_), .A3(new_n684_), .A4(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G43gat), .B1(new_n674_), .B2(new_n443_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT102), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT47), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n711_), .A2(new_n716_), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1330gat));
  NAND2_X1  g517(.A1(new_n684_), .A2(new_n637_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G50gat), .B1(new_n719_), .B2(new_n686_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT103), .Z(new_n721_));
  NAND3_X1  g520(.A1(new_n674_), .A2(new_n471_), .A3(new_n637_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1331gat));
  INV_X1    g522(.A(new_n610_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n653_), .A2(new_n724_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT104), .Z(new_n726_));
  AOI21_X1  g525(.A(new_n631_), .B1(new_n640_), .B2(new_n408_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT105), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n402_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(KEYINPUT105), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n533_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NOR4_X1   g531(.A1(new_n532_), .A2(new_n581_), .A3(new_n631_), .A4(new_n610_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(G57gat), .A3(new_n402_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT106), .Z(G1332gat));
  AOI21_X1  g535(.A(new_n535_), .B1(new_n733_), .B2(new_n658_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n728_), .A2(new_n535_), .A3(new_n658_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1333gat));
  AOI21_X1  g540(.A(new_n547_), .B1(new_n733_), .B2(new_n443_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT109), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n728_), .A2(new_n547_), .A3(new_n443_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1334gat));
  AOI21_X1  g546(.A(new_n256_), .B1(new_n733_), .B2(new_n637_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT50), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n728_), .A2(new_n256_), .A3(new_n637_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1335gat));
  AND3_X1   g550(.A1(new_n727_), .A2(new_n724_), .A3(new_n673_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(new_n455_), .A3(new_n402_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n651_), .B1(new_n640_), .B2(new_n408_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n681_), .B1(new_n680_), .B2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n679_), .B1(new_n754_), .B2(new_n680_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT110), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n677_), .A2(new_n678_), .A3(new_n758_), .A4(new_n681_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n610_), .A2(new_n631_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n581_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n757_), .A2(new_n759_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n757_), .A2(KEYINPUT111), .A3(new_n759_), .A4(new_n762_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n402_), .A3(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n753_), .B1(new_n767_), .B2(new_n455_), .ZN(G1336gat));
  NAND3_X1  g567(.A1(new_n752_), .A2(new_n456_), .A3(new_n658_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n765_), .A2(new_n658_), .A3(new_n766_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n456_), .ZN(G1337gat));
  NAND3_X1  g570(.A1(new_n765_), .A2(new_n443_), .A3(new_n766_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G99gat), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n752_), .A2(new_n443_), .A3(new_n480_), .A4(new_n481_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT51), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(new_n777_), .A3(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n752_), .A2(new_n449_), .A3(new_n637_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT112), .Z(new_n781_));
  NOR2_X1   g580(.A1(new_n761_), .A2(new_n279_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n449_), .B1(new_n682_), .B2(new_n782_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n783_), .A2(KEYINPUT52), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(KEYINPUT52), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g586(.A1(new_n279_), .A2(new_n402_), .A3(new_n363_), .A4(new_n443_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n636_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n591_), .A2(new_n589_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n494_), .A2(new_n584_), .B1(KEYINPUT67), .B2(KEYINPUT12), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n594_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT114), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n592_), .A2(new_n795_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n591_), .A2(new_n589_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n797_), .A2(KEYINPUT55), .A3(new_n588_), .A4(new_n587_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n594_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n794_), .A2(new_n796_), .A3(new_n798_), .A4(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n599_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(KEYINPUT56), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n801_), .B2(new_n802_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n790_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n604_), .A2(new_n606_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n613_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n618_), .A2(new_n620_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n628_), .B1(new_n808_), .B2(new_n623_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n629_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n805_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT57), .B1(new_n812_), .B2(new_n531_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  INV_X1    g613(.A(new_n524_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n529_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n530_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n814_), .B(new_n818_), .C1(new_n805_), .C2(new_n811_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n813_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n810_), .A2(new_n604_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n801_), .A2(new_n802_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n801_), .A2(KEYINPUT56), .A3(new_n802_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n821_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT58), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n810_), .A2(new_n604_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(KEYINPUT115), .A3(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n652_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n580_), .B1(new_n820_), .B2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n651_), .A2(new_n580_), .A3(new_n636_), .A4(new_n610_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n835_), .A2(KEYINPUT113), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT54), .B1(new_n835_), .B2(KEYINPUT113), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n835_), .A2(KEYINPUT113), .A3(new_n839_), .ZN(new_n840_));
  NOR4_X1   g639(.A1(new_n834_), .A2(new_n838_), .A3(KEYINPUT116), .A4(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n631_), .A2(new_n604_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n811_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n531_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n814_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n812_), .A2(KEYINPUT57), .A3(new_n531_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n833_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n840_), .B1(new_n849_), .B2(new_n581_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n838_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n842_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n789_), .B1(new_n841_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT59), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n850_), .A2(new_n851_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n789_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n636_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n853_), .A2(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT117), .B(new_n789_), .C1(new_n841_), .C2(new_n852_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n636_), .A2(G113gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n859_), .B1(new_n863_), .B2(new_n864_), .ZN(G1340gat));
  INV_X1    g664(.A(KEYINPUT60), .ZN(new_n866_));
  AOI21_X1  g665(.A(G120gat), .B1(new_n724_), .B2(new_n866_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT118), .Z(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n866_), .B2(G120gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n861_), .A2(new_n862_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n861_), .A2(KEYINPUT119), .A3(new_n862_), .A4(new_n869_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G120gat), .B1(new_n858_), .B2(new_n610_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT120), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n874_), .A2(new_n878_), .A3(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1341gat));
  OAI21_X1  g679(.A(G127gat), .B1(new_n858_), .B2(new_n581_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n581_), .A2(G127gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n863_), .B2(new_n882_), .ZN(G1342gat));
  OAI21_X1  g682(.A(G134gat), .B1(new_n858_), .B2(new_n651_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n531_), .A2(G134gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n863_), .B2(new_n885_), .ZN(G1343gat));
  INV_X1    g685(.A(new_n852_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n850_), .A2(new_n851_), .A3(new_n842_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n279_), .A2(new_n658_), .A3(new_n409_), .A4(new_n443_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n636_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT121), .B(G141gat), .Z(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1344gat));
  NOR2_X1   g693(.A1(new_n891_), .A2(new_n610_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT122), .B(G148gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1345gat));
  NOR2_X1   g696(.A1(new_n891_), .A2(new_n581_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT61), .B(G155gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n891_), .B2(new_n651_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n531_), .A2(G162gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n891_), .B2(new_n902_), .ZN(G1347gat));
  NAND2_X1  g702(.A1(new_n658_), .A2(new_n403_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n631_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n279_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n907_), .B2(new_n906_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n855_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n286_), .B1(new_n910_), .B2(KEYINPUT124), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(KEYINPUT124), .B2(new_n910_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT62), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n904_), .A2(new_n637_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n855_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n915_), .A2(new_n318_), .A3(new_n631_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n916_), .ZN(G1348gat));
  INV_X1    g716(.A(new_n915_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n287_), .B1(new_n918_), .B2(new_n610_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n637_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n905_), .A2(new_n724_), .A3(G176gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n919_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT125), .ZN(G1349gat));
  NOR3_X1   g723(.A1(new_n918_), .A2(new_n295_), .A3(new_n581_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n920_), .A2(new_n580_), .A3(new_n905_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n281_), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n918_), .B2(new_n651_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n818_), .A2(new_n293_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT126), .Z(new_n930_));
  OAI21_X1  g729(.A(new_n928_), .B1(new_n918_), .B2(new_n930_), .ZN(G1351gat));
  NOR4_X1   g730(.A1(new_n279_), .A2(new_n363_), .A3(new_n402_), .A4(new_n443_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n889_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n631_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n724_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g736(.A1(new_n933_), .A2(new_n580_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  AND2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n938_), .A2(new_n939_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n942_), .A2(KEYINPUT127), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(KEYINPUT127), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n941_), .B1(new_n943_), .B2(new_n944_), .ZN(G1354gat));
  INV_X1    g744(.A(new_n933_), .ZN(new_n946_));
  OAI21_X1  g745(.A(G218gat), .B1(new_n946_), .B2(new_n651_), .ZN(new_n947_));
  OR2_X1    g746(.A1(new_n531_), .A2(G218gat), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n946_), .B2(new_n948_), .ZN(G1355gat));
endmodule


