//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_;
  XNOR2_X1  g000(.A(KEYINPUT18), .B(G64gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT99), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT96), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT22), .B(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT97), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n212_), .B1(new_n215_), .B2(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n217_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n212_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT82), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(G190gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT23), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n223_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n226_), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n229_), .A2(KEYINPUT98), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT98), .B1(new_n229_), .B2(new_n230_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n218_), .B(new_n220_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n222_), .A2(KEYINPUT84), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n222_), .A2(KEYINPUT84), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n227_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n217_), .A2(KEYINPUT24), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  MUX2_X1   g037(.A(new_n237_), .B(KEYINPUT24), .S(new_n238_), .Z(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT25), .B(G183gat), .Z(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT26), .B(G190gat), .Z(new_n241_));
  OAI211_X1 g040(.A(new_n236_), .B(new_n239_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n233_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT91), .B(G197gat), .ZN(new_n244_));
  INV_X1    g043(.A(G204gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G197gat), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n246_), .B(KEYINPUT21), .C1(new_n247_), .C2(new_n245_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(G204gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(G197gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n248_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT21), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n211_), .B1(new_n243_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  AOI211_X1 g058(.A(KEYINPUT99), .B(new_n259_), .C1(new_n233_), .C2(new_n242_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n257_), .B(KEYINPUT93), .ZN(new_n263_));
  INV_X1    g062(.A(G176gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n219_), .B1(new_n213_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT83), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT81), .B(G190gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n236_), .B1(G183gat), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n267_), .B2(KEYINPUT26), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n229_), .B(new_n239_), .C1(new_n271_), .C2(new_n240_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n262_), .B1(new_n263_), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n210_), .B1(new_n261_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT93), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n257_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n269_), .A2(new_n272_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n233_), .A2(new_n259_), .A3(new_n242_), .ZN(new_n280_));
  AND4_X1   g079(.A1(KEYINPUT20), .A2(new_n279_), .A3(new_n210_), .A4(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n207_), .B1(new_n275_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n243_), .A2(new_n257_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT99), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n243_), .A2(new_n211_), .A3(new_n257_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n274_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n281_), .B1(new_n286_), .B2(new_n209_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n207_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT104), .B(KEYINPUT27), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n284_), .A2(new_n210_), .A3(new_n274_), .A4(new_n285_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n279_), .A2(new_n280_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n209_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n207_), .B(KEYINPUT103), .Z(new_n298_));
  AOI22_X1  g097(.A1(new_n287_), .A2(new_n288_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n290_), .A2(new_n292_), .B1(new_n299_), .B2(KEYINPUT27), .ZN(new_n300_));
  NOR3_X1   g099(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT3), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n304_), .B1(new_n305_), .B2(KEYINPUT2), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n305_), .A2(KEYINPUT2), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n305_), .A2(KEYINPUT2), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n303_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n302_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT88), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G155gat), .B(G162gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(KEYINPUT89), .Z(new_n314_));
  NAND4_X1  g113(.A1(new_n302_), .A2(KEYINPUT88), .A3(new_n306_), .A4(new_n309_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n304_), .B1(KEYINPUT1), .B2(new_n317_), .ZN(new_n318_));
  OAI221_X1 g117(.A(new_n318_), .B1(G141gat), .B2(G148gat), .C1(KEYINPUT1), .C2(new_n313_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G127gat), .B(G134gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G113gat), .ZN(new_n322_));
  INV_X1    g121(.A(G120gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT100), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n320_), .A2(new_n325_), .A3(KEYINPUT100), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n326_), .A2(KEYINPUT4), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n330_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(KEYINPUT4), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n333_), .B1(new_n336_), .B2(new_n332_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G85gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(G1gat), .B(G29gat), .Z(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT102), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n333_), .B(new_n341_), .C1(new_n336_), .C2(new_n332_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  OR3_X1    g145(.A1(new_n337_), .A2(new_n344_), .A3(new_n342_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n300_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n320_), .A2(KEYINPUT29), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n257_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(G228gat), .A3(G233gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(G78gat), .B(G106gat), .Z(new_n353_));
  NAND2_X1  g152(.A1(G228gat), .A2(G233gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n277_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n353_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n359_));
  OR3_X1    g158(.A1(new_n320_), .A2(KEYINPUT29), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G22gat), .B(G50gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n359_), .B1(new_n320_), .B2(KEYINPUT29), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT94), .B1(new_n358_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G15gat), .B(G43gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n278_), .A2(KEYINPUT30), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n278_), .A2(KEYINPUT30), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n278_), .A2(KEYINPUT30), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n373_), .B1(new_n376_), .B2(new_n370_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n369_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n324_), .B(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n374_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n370_), .A3(new_n373_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n369_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n378_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n380_), .B1(new_n378_), .B2(new_n384_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT95), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n388_), .B1(new_n357_), .B2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n352_), .A2(KEYINPUT95), .A3(new_n355_), .A4(new_n353_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n365_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT94), .ZN(new_n393_));
  OAI221_X1 g192(.A(new_n393_), .B1(new_n363_), .B2(new_n364_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n394_));
  AND4_X1   g193(.A1(new_n366_), .A2(new_n387_), .A3(new_n392_), .A4(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT105), .B1(new_n349_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT105), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n395_), .A2(new_n300_), .A3(new_n348_), .A4(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n366_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n349_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n290_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n342_), .B1(new_n336_), .B2(new_n332_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n332_), .B2(new_n331_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n343_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n337_), .A2(KEYINPUT33), .A3(new_n342_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n403_), .A2(new_n405_), .A3(new_n407_), .A4(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n288_), .A2(KEYINPUT32), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n297_), .A2(new_n410_), .ZN(new_n411_));
  OR3_X1    g210(.A1(new_n275_), .A2(new_n410_), .A3(new_n281_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n346_), .A2(new_n347_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n401_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n409_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n387_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n402_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n400_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT74), .B(G43gat), .ZN(new_n419_));
  INV_X1    g218(.A(G50gat), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n419_), .A2(new_n420_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G29gat), .B(G36gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT78), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G15gat), .B(G22gat), .ZN(new_n427_));
  INV_X1    g226(.A(G1gat), .ZN(new_n428_));
  INV_X1    g227(.A(G8gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT14), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G1gat), .B(G8gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n431_), .B(new_n432_), .Z(new_n433_));
  XNOR2_X1  g232(.A(new_n426_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G229gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n426_), .A2(new_n433_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n425_), .B(KEYINPUT15), .ZN(new_n439_));
  INV_X1    g238(.A(new_n433_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n438_), .A2(new_n441_), .A3(new_n435_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G113gat), .B(G141gat), .ZN(new_n444_));
  INV_X1    g243(.A(G169gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(new_n247_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(KEYINPUT79), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT80), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n443_), .B(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT10), .B(G99gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT64), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT65), .B1(new_n454_), .B2(G106gat), .ZN(new_n455_));
  INV_X1    g254(.A(G85gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT66), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT9), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(G92gat), .ZN(new_n459_));
  INV_X1    g258(.A(G92gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT66), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n456_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G85gat), .B(G92gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI211_X1 g269(.A(new_n462_), .B(new_n468_), .C1(KEYINPUT9), .C2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT64), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n453_), .B(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT65), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n455_), .A2(new_n471_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT67), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n467_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n464_), .A2(new_n466_), .A3(KEYINPUT67), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n481_));
  INV_X1    g280(.A(G99gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n475_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n483_), .A2(KEYINPUT68), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT68), .B1(new_n483_), .B2(new_n484_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n479_), .B(new_n480_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n470_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT69), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT69), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n487_), .A2(new_n490_), .A3(new_n470_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(KEYINPUT8), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n484_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT8), .B1(new_n495_), .B2(new_n467_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n470_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n477_), .B1(new_n492_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n502_));
  XOR2_X1   g301(.A(G71gat), .B(G78gat), .Z(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n502_), .A2(new_n503_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n498_), .A2(new_n499_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT70), .ZN(new_n508_));
  INV_X1    g307(.A(new_n497_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n464_), .A2(new_n466_), .A3(KEYINPUT67), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT67), .B1(new_n464_), .B2(new_n466_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT68), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n483_), .A2(KEYINPUT68), .A3(new_n484_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI211_X1 g315(.A(KEYINPUT69), .B(new_n469_), .C1(new_n512_), .C2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n490_), .B1(new_n487_), .B2(new_n470_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n509_), .B1(new_n519_), .B2(KEYINPUT8), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n508_), .B1(new_n520_), .B2(new_n477_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n506_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n498_), .A2(KEYINPUT70), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n507_), .B1(new_n524_), .B2(new_n499_), .ZN(new_n525_));
  AND2_X1   g324(.A1(G230gat), .A2(G233gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n521_), .A2(new_n523_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n527_), .B2(new_n506_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n522_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n526_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G120gat), .B(G148gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  NAND3_X1  g336(.A1(new_n529_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT72), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n529_), .A2(new_n532_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n537_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n541_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(KEYINPUT72), .A3(new_n538_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT13), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(KEYINPUT73), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n452_), .B1(new_n548_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n418_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n527_), .A2(new_n425_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT34), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT35), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n439_), .B1(new_n520_), .B2(new_n477_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(KEYINPUT35), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n562_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT75), .B(G134gat), .ZN(new_n565_));
  INV_X1    g364(.A(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT36), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n563_), .A2(new_n564_), .A3(new_n571_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n563_), .A2(new_n564_), .B1(new_n570_), .B2(new_n569_), .ZN(new_n573_));
  OAI211_X1 g372(.A(KEYINPUT76), .B(KEYINPUT37), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n563_), .A2(new_n564_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n569_), .A2(new_n570_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n563_), .A2(new_n564_), .A3(new_n571_), .ZN(new_n578_));
  OR2_X1    g377(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n579_));
  NAND2_X1  g378(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .A4(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n433_), .B(new_n506_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT16), .B(G183gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G211gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n589_), .B(new_n590_), .Z(new_n591_));
  OAI21_X1  g390(.A(new_n586_), .B1(new_n587_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(KEYINPUT17), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n592_), .B1(new_n586_), .B2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT77), .Z(new_n595_));
  NOR2_X1   g394(.A1(new_n583_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n555_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n348_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n428_), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT38), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n572_), .A2(new_n573_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n554_), .A2(new_n595_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G1gat), .B1(new_n605_), .B2(new_n348_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT106), .ZN(G1324gat));
  INV_X1    g407(.A(new_n300_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n604_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(G8gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT39), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n598_), .A2(new_n429_), .A3(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(G1325gat));
  OAI21_X1  g415(.A(G15gat), .B1(new_n605_), .B2(new_n416_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT41), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n597_), .A2(G15gat), .A3(new_n416_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1326gat));
  INV_X1    g419(.A(G22gat), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n604_), .B2(new_n401_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT42), .Z(new_n623_));
  NAND2_X1  g422(.A1(new_n401_), .A2(new_n621_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT107), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n623_), .B1(new_n597_), .B2(new_n625_), .ZN(G1327gat));
  INV_X1    g425(.A(KEYINPUT44), .ZN(new_n627_));
  INV_X1    g426(.A(new_n595_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n553_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n387_), .B1(new_n349_), .B2(new_n401_), .ZN(new_n630_));
  AOI22_X1  g429(.A1(new_n397_), .A2(new_n399_), .B1(new_n630_), .B2(new_n415_), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT43), .B1(new_n631_), .B2(new_n582_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n418_), .A2(new_n633_), .A3(new_n583_), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n628_), .B(new_n629_), .C1(new_n632_), .C2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT108), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n627_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n634_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n595_), .A3(new_n553_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n348_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(G29gat), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n554_), .A2(new_n628_), .A3(new_n602_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n599_), .A2(new_n642_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT109), .Z(new_n646_));
  OAI22_X1  g445(.A1(new_n641_), .A2(new_n642_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT110), .ZN(G1328gat));
  INV_X1    g447(.A(KEYINPUT112), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n649_), .A2(KEYINPUT46), .ZN(new_n650_));
  INV_X1    g449(.A(G36gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n643_), .A2(new_n651_), .A3(new_n609_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT45), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n300_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n650_), .B(new_n653_), .C1(new_n654_), .C2(new_n651_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT111), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n649_), .B1(new_n656_), .B2(KEYINPUT46), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n655_), .B(new_n657_), .ZN(G1329gat));
  INV_X1    g457(.A(KEYINPUT47), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n637_), .A2(new_n640_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n387_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G43gat), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n644_), .A2(G43gat), .A3(new_n416_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n659_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT47), .B(new_n663_), .C1(new_n661_), .C2(G43gat), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1330gat));
  NAND3_X1  g466(.A1(new_n643_), .A2(new_n420_), .A3(new_n401_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n414_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(new_n420_), .ZN(G1331gat));
  NAND2_X1  g469(.A1(new_n548_), .A2(new_n552_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n451_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n672_), .A2(new_n628_), .A3(new_n602_), .A4(new_n418_), .ZN(new_n673_));
  INV_X1    g472(.A(G57gat), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n348_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n418_), .A2(new_n452_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT113), .ZN(new_n677_));
  INV_X1    g476(.A(new_n671_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n677_), .A2(new_n678_), .A3(new_n596_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n599_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n675_), .B1(new_n680_), .B2(new_n674_), .ZN(G1332gat));
  OAI21_X1  g480(.A(G64gat), .B1(new_n673_), .B2(new_n300_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT114), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT48), .ZN(new_n684_));
  INV_X1    g483(.A(G64gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n679_), .A2(new_n685_), .A3(new_n609_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1333gat));
  NOR2_X1   g486(.A1(new_n416_), .A2(G71gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT115), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n679_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G71gat), .B1(new_n673_), .B2(new_n416_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT49), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1334gat));
  INV_X1    g492(.A(G78gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n679_), .A2(new_n694_), .A3(new_n401_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G78gat), .B1(new_n673_), .B2(new_n414_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT50), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1335gat));
  NOR2_X1   g497(.A1(new_n602_), .A2(new_n628_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n677_), .A2(new_n678_), .A3(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(new_n456_), .A3(new_n599_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n638_), .A2(new_n595_), .A3(new_n672_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT116), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n703_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT117), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(KEYINPUT117), .A3(new_n705_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n348_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n701_), .B1(new_n710_), .B2(new_n456_), .ZN(G1336gat));
  AOI21_X1  g510(.A(G92gat), .B1(new_n700_), .B2(new_n609_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n457_), .A2(G92gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n461_), .B1(new_n300_), .B2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n712_), .B1(new_n713_), .B2(new_n715_), .ZN(G1337gat));
  NAND3_X1  g515(.A1(new_n704_), .A2(new_n387_), .A3(new_n705_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G99gat), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n677_), .A2(new_n473_), .A3(new_n678_), .A4(new_n699_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT118), .B1(new_n719_), .B2(new_n416_), .ZN(new_n720_));
  OR3_X1    g519(.A1(new_n719_), .A2(KEYINPUT118), .A3(new_n416_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n718_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT51), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n718_), .A2(new_n724_), .A3(new_n720_), .A4(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1338gat));
  NAND3_X1  g525(.A1(new_n700_), .A2(new_n475_), .A3(new_n401_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n702_), .A2(new_n414_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(G106gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G106gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT53), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n734_), .B(new_n727_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1339gat));
  NOR2_X1   g535(.A1(new_n595_), .A2(new_n451_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT119), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n582_), .B(new_n739_), .C1(new_n547_), .C2(new_n551_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT54), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n527_), .A2(new_n506_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n507_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n743_), .B(new_n744_), .C1(new_n530_), .C2(KEYINPUT12), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n526_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n525_), .A2(new_n747_), .A3(new_n528_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT120), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT120), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n746_), .B(new_n752_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n751_), .A2(new_n541_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n541_), .A4(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n434_), .A2(new_n436_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n438_), .A2(new_n441_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT121), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n759_), .B1(new_n762_), .B2(new_n436_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(new_n448_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n538_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n443_), .A2(new_n447_), .ZN(new_n766_));
  OR3_X1    g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n758_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n758_), .A2(KEYINPUT58), .A3(new_n768_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n583_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n451_), .A2(new_n538_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n764_), .A2(new_n766_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n545_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n602_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT57), .B(new_n602_), .C1(new_n775_), .C2(new_n777_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n773_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n742_), .B1(new_n782_), .B2(new_n595_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n609_), .A2(new_n348_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n785_), .A2(new_n396_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n783_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G113gat), .B1(new_n788_), .B2(new_n451_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n780_), .A2(new_n781_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT58), .B1(new_n758_), .B2(new_n768_), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n770_), .B(new_n767_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n582_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n595_), .B1(new_n790_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n742_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(KEYINPUT59), .A3(new_n786_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n783_), .B2(new_n787_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n452_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n789_), .B1(new_n800_), .B2(G113gat), .ZN(G1340gat));
  AOI21_X1  g600(.A(KEYINPUT59), .B1(new_n796_), .B2(new_n786_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n783_), .A2(new_n798_), .A3(new_n787_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n678_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT122), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT122), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(new_n678_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(G120gat), .A3(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n323_), .B1(new_n671_), .B2(KEYINPUT60), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n788_), .B(new_n809_), .C1(KEYINPUT60), .C2(new_n323_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1341gat));
  AOI21_X1  g610(.A(G127gat), .B1(new_n788_), .B2(new_n628_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n595_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g613(.A(G134gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n788_), .A2(new_n815_), .A3(new_n603_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n582_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n815_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT123), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT123), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n816_), .B(new_n820_), .C1(new_n817_), .C2(new_n815_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1343gat));
  NOR3_X1   g621(.A1(new_n783_), .A2(new_n414_), .A3(new_n387_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n451_), .A3(new_n784_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT124), .B(G141gat), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(G1344gat));
  NAND3_X1  g625(.A1(new_n823_), .A2(new_n678_), .A3(new_n784_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g627(.A1(new_n823_), .A2(new_n628_), .A3(new_n784_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1346gat));
  AND2_X1   g630(.A1(new_n823_), .A2(new_n784_), .ZN(new_n832_));
  AOI21_X1  g631(.A(G162gat), .B1(new_n832_), .B2(new_n603_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n582_), .A2(new_n566_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(new_n834_), .ZN(G1347gat));
  NOR2_X1   g634(.A1(new_n599_), .A2(new_n300_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n395_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n783_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n445_), .B1(new_n838_), .B2(new_n451_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n840_), .ZN(new_n842_));
  OR3_X1    g641(.A1(new_n783_), .A2(KEYINPUT125), .A3(new_n837_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT125), .B1(new_n783_), .B2(new_n837_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n452_), .A2(new_n215_), .ZN(new_n846_));
  OAI22_X1  g645(.A1(new_n841_), .A2(new_n842_), .B1(new_n845_), .B2(new_n846_), .ZN(G1348gat));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n844_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(new_n264_), .A3(new_n678_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n783_), .A2(new_n671_), .A3(new_n837_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n264_), .B2(new_n850_), .ZN(G1349gat));
  AND2_X1   g650(.A1(new_n628_), .A2(new_n240_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n848_), .A2(KEYINPUT126), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT126), .B1(new_n848_), .B2(new_n852_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G183gat), .B1(new_n838_), .B2(new_n628_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(G1350gat));
  OAI21_X1  g655(.A(G190gat), .B1(new_n845_), .B2(new_n582_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n602_), .A2(new_n241_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n845_), .B2(new_n858_), .ZN(G1351gat));
  NAND3_X1  g658(.A1(new_n823_), .A2(new_n451_), .A3(new_n836_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g660(.A1(new_n823_), .A2(new_n678_), .A3(new_n836_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g662(.A1(new_n823_), .A2(new_n836_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n628_), .A3(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT127), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n866_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n864_), .A2(new_n628_), .A3(new_n868_), .A4(new_n865_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1354gat));
  AOI21_X1  g671(.A(G218gat), .B1(new_n864_), .B2(new_n603_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n583_), .A2(G218gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n864_), .B2(new_n874_), .ZN(G1355gat));
endmodule


