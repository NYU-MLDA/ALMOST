//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n569_,
    new_n570_, new_n571_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n795_, new_n796_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_;
  INV_X1    g000(.A(KEYINPUT104), .ZN(new_n202_));
  OR2_X1    g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  AND3_X1   g003(.A1(new_n203_), .A2(KEYINPUT24), .A3(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n203_), .A2(KEYINPUT24), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT25), .B(G183gat), .Z(new_n212_));
  OAI211_X1 g011(.A(new_n207_), .B(new_n209_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(G183gat), .B2(G190gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT22), .B(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n204_), .B(KEYINPUT93), .Z(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n213_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G197gat), .B(G204gat), .Z(new_n222_));
  INV_X1    g021(.A(KEYINPUT90), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT21), .ZN(new_n224_));
  XOR2_X1   g023(.A(G211gat), .B(G218gat), .Z(new_n225_));
  OAI22_X1  g024(.A1(new_n224_), .A2(new_n225_), .B1(KEYINPUT21), .B2(new_n222_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n224_), .A2(new_n225_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT94), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n218_), .A2(new_n204_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT83), .B(G183gat), .ZN(new_n232_));
  INV_X1    g031(.A(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n231_), .A2(KEYINPUT84), .B1(new_n234_), .B2(new_n214_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(KEYINPUT84), .B2(new_n231_), .ZN(new_n236_));
  MUX2_X1   g035(.A(G183gat), .B(new_n232_), .S(KEYINPUT25), .Z(new_n237_));
  OAI211_X1 g036(.A(new_n209_), .B(new_n207_), .C1(new_n237_), .C2(new_n211_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n230_), .B(KEYINPUT20), .C1(new_n239_), .C2(new_n228_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n241_));
  NAND2_X1  g040(.A1(G226gat), .A2(G233gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT20), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n221_), .A2(new_n228_), .ZN(new_n246_));
  AOI211_X1 g045(.A(new_n245_), .B(new_n243_), .C1(new_n246_), .C2(KEYINPUT95), .ZN(new_n247_));
  INV_X1    g046(.A(new_n228_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(new_n238_), .B2(new_n236_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n247_), .B(new_n250_), .C1(KEYINPUT95), .C2(new_n246_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n244_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT18), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G64gat), .B(G92gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n254_), .B(new_n255_), .Z(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n252_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n244_), .A2(new_n256_), .A3(new_n251_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n202_), .B1(new_n261_), .B2(KEYINPUT27), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT27), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(KEYINPUT104), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n246_), .A2(KEYINPUT20), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n243_), .B1(new_n266_), .B2(new_n249_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n267_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n257_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(KEYINPUT27), .A3(new_n259_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n273_));
  INV_X1    g072(.A(G99gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G227gat), .A2(G233gat), .ZN(new_n276_));
  INV_X1    g075(.A(G15gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G71gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n275_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G127gat), .B(G134gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT87), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G113gat), .B(G120gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n282_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n280_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT85), .B(G43gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT86), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT31), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n286_), .B(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G141gat), .B(G148gat), .Z(new_n291_));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT1), .ZN(new_n293_));
  OR2_X1    g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n292_), .A2(KEYINPUT1), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n291_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n297_), .B(KEYINPUT88), .Z(new_n298_));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(KEYINPUT3), .Z(new_n300_));
  NAND2_X1  g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n301_), .B(KEYINPUT2), .Z(new_n302_));
  OAI211_X1 g101(.A(new_n292_), .B(new_n294_), .C1(new_n300_), .C2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n248_), .B1(new_n304_), .B2(KEYINPUT29), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G228gat), .A2(G233gat), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n306_), .A2(KEYINPUT91), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n305_), .A2(G78gat), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(G78gat), .B1(new_n305_), .B2(new_n307_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n309_), .A2(G106gat), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(G106gat), .B1(new_n309_), .B2(new_n310_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n304_), .A2(KEYINPUT29), .ZN(new_n313_));
  XOR2_X1   g112(.A(G22gat), .B(G50gat), .Z(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  OR3_X1    g114(.A1(new_n311_), .A2(new_n312_), .A3(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n306_), .A2(KEYINPUT91), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n315_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n316_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n319_), .B1(new_n316_), .B2(new_n320_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n304_), .A2(new_n285_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(KEYINPUT4), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n298_), .A2(new_n303_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n285_), .A2(KEYINPUT96), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n282_), .B(new_n283_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT96), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n327_), .A2(new_n328_), .A3(new_n331_), .A4(KEYINPUT97), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n327_), .A2(new_n328_), .A3(new_n331_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT97), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n325_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n332_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n326_), .B1(new_n336_), .B2(KEYINPUT4), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G225gat), .A2(G233gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(KEYINPUT98), .Z(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT99), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G85gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT0), .B(G57gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  NAND2_X1  g144(.A1(new_n336_), .A2(new_n338_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n336_), .A2(KEYINPUT4), .ZN(new_n347_));
  INV_X1    g146(.A(new_n326_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n347_), .A2(KEYINPUT99), .A3(new_n348_), .A4(new_n339_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n341_), .A2(new_n345_), .A3(new_n346_), .A4(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT103), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n346_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n345_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n340_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT103), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n353_), .B2(new_n340_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n352_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n272_), .A2(new_n290_), .A3(new_n324_), .A4(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n323_), .A2(new_n352_), .A3(new_n357_), .A4(new_n356_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n361_), .A2(new_n271_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT100), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT33), .B1(new_n355_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT33), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n350_), .A2(KEYINPUT100), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n337_), .A2(new_n338_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n345_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n260_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT101), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT101), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n364_), .A2(new_n366_), .A3(new_n372_), .A4(new_n369_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n256_), .A2(KEYINPUT32), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n244_), .A2(new_n251_), .A3(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(KEYINPUT102), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n375_), .A2(KEYINPUT102), .ZN(new_n377_));
  INV_X1    g176(.A(new_n374_), .ZN(new_n378_));
  AOI211_X1 g177(.A(new_n376_), .B(new_n377_), .C1(new_n378_), .C2(new_n268_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n358_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n371_), .A2(new_n373_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n362_), .B1(new_n381_), .B2(new_n324_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n360_), .B1(new_n382_), .B2(new_n290_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT80), .B(G1gat), .ZN(new_n384_));
  INV_X1    g183(.A(G8gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT14), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G15gat), .B(G22gat), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G8gat), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n389_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G43gat), .B(G50gat), .Z(new_n393_));
  XNOR2_X1  g192(.A(G29gat), .B(G36gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n392_), .B(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G229gat), .A2(G233gat), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n392_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n399_), .A2(new_n395_), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n395_), .B(KEYINPUT15), .Z(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n397_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n398_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G113gat), .B(G141gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G169gat), .B(G197gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n404_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n383_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G57gat), .B(G64gat), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n413_), .A2(KEYINPUT11), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(KEYINPUT11), .ZN(new_n415_));
  XOR2_X1   g214(.A(G71gat), .B(G78gat), .Z(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n415_), .A2(new_n416_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT65), .B(G92gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G85gat), .ZN(new_n422_));
  OR3_X1    g221(.A1(new_n421_), .A2(KEYINPUT9), .A3(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G85gat), .B(G92gat), .Z(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT9), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT64), .B(G106gat), .Z(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT10), .B(G99gat), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G99gat), .A2(G106gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT6), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n423_), .A2(new_n425_), .A3(new_n428_), .A4(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT7), .ZN(new_n432_));
  INV_X1    g231(.A(G106gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n274_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT67), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT67), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n436_), .A2(new_n432_), .A3(new_n274_), .A4(new_n433_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT66), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT66), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n441_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(new_n430_), .A3(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n445_));
  AND2_X1   g244(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n444_), .B(new_n424_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT8), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT69), .B(KEYINPUT6), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n429_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n429_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n452_), .A2(KEYINPUT69), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(KEYINPUT69), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n451_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n438_), .A2(new_n443_), .A3(new_n450_), .A4(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n448_), .B1(new_n456_), .B2(new_n424_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT70), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n447_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  AOI211_X1 g258(.A(KEYINPUT70), .B(new_n448_), .C1(new_n456_), .C2(new_n424_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n419_), .B(new_n431_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G230gat), .A2(G233gat), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n431_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT12), .ZN(new_n465_));
  INV_X1    g264(.A(new_n419_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n463_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT72), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n464_), .A2(new_n466_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT71), .ZN(new_n473_));
  INV_X1    g272(.A(new_n462_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT71), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n461_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n473_), .B(new_n474_), .C1(new_n472_), .C2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT72), .B(new_n463_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n471_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G120gat), .B(G148gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT5), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G176gat), .B(G204gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n479_), .A2(KEYINPUT73), .A3(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n471_), .A2(new_n477_), .A3(new_n478_), .A4(new_n484_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT73), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n489_), .B1(new_n479_), .B2(new_n484_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n491_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G231gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n419_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(new_n399_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G127gat), .B(G155gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT16), .ZN(new_n501_));
  XOR2_X1   g300(.A(G183gat), .B(G211gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n498_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(KEYINPUT17), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT34), .Z(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT74), .B(KEYINPUT35), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n464_), .A2(new_n395_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n464_), .A2(new_n401_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n509_), .A2(new_n510_), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n514_), .B(KEYINPUT75), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT77), .ZN(new_n516_));
  AND4_X1   g315(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .A4(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n511_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT76), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT76), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n512_), .A2(new_n520_), .A3(new_n511_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n521_), .A3(new_n513_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n517_), .B1(new_n522_), .B2(new_n515_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G190gat), .B(G218gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G134gat), .B(G162gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(KEYINPUT36), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n526_), .B(KEYINPUT36), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT79), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n523_), .B2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT78), .B1(new_n523_), .B2(new_n530_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT37), .A3(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n523_), .A2(new_n530_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n534_), .B(new_n528_), .C1(KEYINPUT78), .C2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n507_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n495_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT81), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n412_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n358_), .A2(KEYINPUT105), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n358_), .A2(KEYINPUT105), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n384_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT38), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT106), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n531_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n534_), .A2(KEYINPUT106), .A3(new_n528_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n383_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n495_), .A2(new_n411_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(new_n507_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(G1gat), .B1(new_n557_), .B2(new_n359_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n546_), .A2(new_n547_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n548_), .A2(new_n558_), .A3(new_n559_), .ZN(G1324gat));
  NAND3_X1  g359(.A1(new_n541_), .A2(new_n385_), .A3(new_n271_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n554_), .A2(new_n556_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n271_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n563_), .A2(G8gat), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n563_), .B2(G8gat), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n561_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g367(.A(new_n277_), .B1(new_n562_), .B2(new_n290_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT41), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n541_), .A2(new_n277_), .A3(new_n290_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(G1326gat));
  OAI21_X1  g371(.A(G22gat), .B1(new_n557_), .B2(new_n324_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT42), .ZN(new_n574_));
  OR3_X1    g373(.A1(new_n540_), .A2(G22gat), .A3(new_n324_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT108), .ZN(G1327gat));
  NOR2_X1   g376(.A1(new_n555_), .A2(new_n506_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT43), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n533_), .A2(new_n536_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n383_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n579_), .B1(new_n383_), .B2(new_n581_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n578_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT44), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(KEYINPUT44), .B(new_n578_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G29gat), .B1(new_n588_), .B2(new_n544_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n552_), .A2(new_n507_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT109), .Z(new_n591_));
  NAND3_X1  g390(.A1(new_n412_), .A2(new_n495_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT110), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n412_), .A2(KEYINPUT110), .A3(new_n495_), .A4(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n359_), .A2(G29gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT111), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n589_), .B1(new_n596_), .B2(new_n598_), .ZN(G1328gat));
  NOR2_X1   g398(.A1(new_n272_), .A2(G36gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n594_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G36gat), .B1(new_n588_), .B2(new_n272_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT46), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(new_n604_), .A3(KEYINPUT46), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1329gat));
  NAND4_X1  g408(.A1(new_n586_), .A2(G43gat), .A3(new_n290_), .A4(new_n587_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n594_), .A2(new_n290_), .A3(new_n595_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT113), .ZN(new_n612_));
  INV_X1    g411(.A(G43gat), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n612_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n610_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT47), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT47), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n618_), .B(new_n610_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(G1330gat));
  INV_X1    g419(.A(G50gat), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n588_), .A2(new_n621_), .A3(new_n324_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n594_), .A2(new_n323_), .A3(new_n595_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n621_), .B2(new_n623_), .ZN(G1331gat));
  NOR2_X1   g423(.A1(new_n495_), .A2(new_n411_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n554_), .A2(new_n506_), .A3(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G57gat), .B1(new_n626_), .B2(new_n359_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n383_), .A2(new_n625_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n537_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n544_), .A2(G57gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n627_), .B1(new_n629_), .B2(new_n630_), .ZN(G1332gat));
  OAI21_X1  g430(.A(G64gat), .B1(new_n626_), .B2(new_n272_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT48), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n272_), .A2(G64gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n633_), .B1(new_n629_), .B2(new_n634_), .ZN(G1333gat));
  INV_X1    g434(.A(new_n290_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G71gat), .B1(new_n626_), .B2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n636_), .A2(G71gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n639_), .B1(new_n629_), .B2(new_n640_), .ZN(G1334gat));
  OAI21_X1  g440(.A(G78gat), .B1(new_n626_), .B2(new_n324_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n324_), .A2(G78gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n629_), .B2(new_n645_), .ZN(G1335gat));
  NAND2_X1  g445(.A1(new_n625_), .A2(new_n507_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n383_), .A2(new_n581_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT43), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n383_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n647_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n422_), .B1(new_n651_), .B2(new_n358_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n628_), .A2(new_n591_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(G85gat), .A3(new_n544_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n652_), .A2(new_n654_), .ZN(G1336gat));
  INV_X1    g454(.A(new_n653_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G92gat), .B1(new_n656_), .B2(new_n271_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n272_), .A2(new_n421_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n651_), .B2(new_n658_), .ZN(G1337gat));
  AOI21_X1  g458(.A(new_n274_), .B1(new_n651_), .B2(new_n290_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n653_), .A2(new_n636_), .A3(new_n427_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT116), .ZN(new_n662_));
  OAI22_X1  g461(.A1(new_n660_), .A2(new_n661_), .B1(new_n662_), .B2(KEYINPUT51), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(KEYINPUT51), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(G1338gat));
  INV_X1    g464(.A(new_n647_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n323_), .B(new_n666_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT117), .ZN(new_n668_));
  OAI21_X1  g467(.A(G106gat), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT117), .B1(new_n651_), .B2(new_n323_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT52), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n651_), .A2(KEYINPUT117), .A3(new_n323_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n667_), .A2(new_n668_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT52), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .A4(G106gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n653_), .A2(new_n324_), .A3(new_n426_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT53), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT53), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n676_), .A2(new_n680_), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1339gat));
  NOR3_X1   g481(.A1(new_n636_), .A2(new_n323_), .A3(new_n271_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n545_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT121), .ZN(new_n685_));
  INV_X1    g484(.A(new_n397_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n400_), .A2(new_n686_), .A3(new_n402_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n396_), .A2(new_n686_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n407_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n404_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(new_n407_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n490_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n489_), .A2(new_n411_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT55), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n471_), .A2(new_n694_), .A3(new_n478_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT118), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n471_), .A2(KEYINPUT118), .A3(new_n694_), .A4(new_n478_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n469_), .A2(new_n694_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n461_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n462_), .B1(new_n700_), .B2(KEYINPUT119), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT119), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n702_), .B(new_n461_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n699_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n697_), .A2(new_n698_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n483_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT56), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n705_), .A2(KEYINPUT56), .A3(new_n483_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n693_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n692_), .B1(new_n710_), .B2(KEYINPUT120), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n410_), .B1(new_n485_), .B2(new_n488_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n705_), .A2(KEYINPUT56), .A3(new_n483_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT56), .B1(new_n705_), .B2(new_n483_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT120), .B(new_n712_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n553_), .B1(new_n711_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT57), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT120), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(new_n715_), .A3(new_n692_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n552_), .A2(new_n718_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n489_), .A2(new_n691_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n725_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT58), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n580_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n725_), .B(KEYINPUT58), .C1(new_n714_), .C2(new_n713_), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n723_), .A2(new_n724_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n506_), .B1(new_n719_), .B2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n537_), .A2(new_n492_), .A3(new_n410_), .A4(new_n493_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT54), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n685_), .B1(new_n731_), .B2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n724_), .B1(new_n711_), .B2(new_n716_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n728_), .A2(new_n729_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT57), .B1(new_n723_), .B2(new_n553_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n507_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(KEYINPUT121), .A3(new_n733_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n684_), .B1(new_n735_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G113gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n743_), .A3(new_n411_), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT59), .B(new_n684_), .C1(new_n740_), .C2(new_n733_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n684_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n731_), .A2(new_n734_), .A3(new_n685_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT121), .B1(new_n740_), .B2(new_n733_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(KEYINPUT122), .A3(KEYINPUT59), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT122), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT59), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n742_), .B2(new_n752_), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n410_), .B(new_n745_), .C1(new_n750_), .C2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n744_), .B1(new_n754_), .B2(new_n743_), .ZN(G1340gat));
  INV_X1    g554(.A(KEYINPUT123), .ZN(new_n756_));
  INV_X1    g555(.A(G120gat), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n750_), .A2(new_n753_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n745_), .A2(new_n495_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n757_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT60), .ZN(new_n761_));
  AOI21_X1  g560(.A(G120gat), .B1(new_n494_), .B2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n761_), .B2(G120gat), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n742_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n756_), .B1(new_n760_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n759_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT123), .B(new_n764_), .C1(new_n768_), .C2(new_n757_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(G1341gat));
  INV_X1    g569(.A(G127gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n742_), .A2(new_n771_), .A3(new_n506_), .ZN(new_n772_));
  AOI211_X1 g571(.A(new_n507_), .B(new_n745_), .C1(new_n750_), .C2(new_n753_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(new_n771_), .ZN(G1342gat));
  NAND2_X1  g573(.A1(new_n581_), .A2(G134gat), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT124), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI211_X1 g576(.A(new_n745_), .B(new_n777_), .C1(new_n750_), .C2(new_n753_), .ZN(new_n778_));
  AOI21_X1  g577(.A(G134gat), .B1(new_n742_), .B2(new_n552_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT125), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n745_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n758_), .A2(new_n781_), .A3(new_n776_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT125), .ZN(new_n783_));
  INV_X1    g582(.A(new_n779_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n780_), .A2(new_n785_), .ZN(G1343gat));
  AOI21_X1  g585(.A(new_n290_), .B1(new_n735_), .B2(new_n741_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n544_), .A2(new_n324_), .A3(new_n271_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n411_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n494_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g593(.A1(new_n789_), .A2(new_n507_), .ZN(new_n795_));
  XOR2_X1   g594(.A(KEYINPUT61), .B(G155gat), .Z(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(G1346gat));
  OAI21_X1  g596(.A(G162gat), .B1(new_n789_), .B2(new_n580_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n553_), .A2(G162gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n789_), .B2(new_n799_), .ZN(G1347gat));
  NAND2_X1  g599(.A1(new_n740_), .A2(new_n733_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n545_), .A2(new_n636_), .A3(new_n272_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(new_n324_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n411_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n806_));
  INV_X1    g605(.A(new_n216_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n805_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT62), .B1(new_n805_), .B2(G169gat), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1348gat));
  AOI21_X1  g609(.A(G176gat), .B1(new_n804_), .B2(new_n494_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n323_), .B1(new_n735_), .B2(new_n741_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n802_), .A2(G176gat), .A3(new_n494_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n811_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT126), .Z(G1349gat));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n506_), .A3(new_n802_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n506_), .A2(new_n212_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n817_), .A2(new_n232_), .B1(new_n804_), .B2(new_n818_), .ZN(G1350gat));
  INV_X1    g618(.A(new_n804_), .ZN(new_n820_));
  OAI21_X1  g619(.A(G190gat), .B1(new_n820_), .B2(new_n580_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n552_), .A2(new_n210_), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n822_), .B(KEYINPUT127), .Z(new_n823_));
  OAI21_X1  g622(.A(new_n821_), .B1(new_n820_), .B2(new_n823_), .ZN(G1351gat));
  NOR2_X1   g623(.A1(new_n272_), .A2(new_n361_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n787_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n411_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n494_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g630(.A1(new_n826_), .A2(new_n507_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n832_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT63), .B(G211gat), .Z(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(new_n834_), .ZN(G1354gat));
  OAI21_X1  g634(.A(G218gat), .B1(new_n826_), .B2(new_n580_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n553_), .A2(G218gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n826_), .B2(new_n837_), .ZN(G1355gat));
endmodule


