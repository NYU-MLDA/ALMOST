//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n908_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_;
  INV_X1    g000(.A(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT6), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT10), .B(G99gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT64), .ZN(new_n210_));
  OR2_X1    g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT9), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  OAI221_X1 g013(.A(new_n207_), .B1(G106gat), .B2(new_n208_), .C1(new_n210_), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT8), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR3_X1   g017(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT65), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n202_), .A3(new_n203_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n217_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n207_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n211_), .A2(new_n213_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n216_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(new_n217_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI211_X1 g029(.A(KEYINPUT8), .B(new_n226_), .C1(new_n230_), .C2(new_n207_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n215_), .B1(new_n228_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT66), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G57gat), .B(G64gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT11), .ZN(new_n235_));
  XOR2_X1   g034(.A(G71gat), .B(G78gat), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n234_), .A2(KEYINPUT11), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n235_), .A2(new_n236_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n242_), .B(new_n215_), .C1(new_n228_), .C2(new_n231_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n233_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT12), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n228_), .B2(new_n231_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n230_), .A2(new_n207_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n216_), .A3(new_n227_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n229_), .A2(KEYINPUT65), .B1(new_n204_), .B2(new_n206_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n226_), .B1(new_n251_), .B2(new_n224_), .ZN(new_n252_));
  OAI211_X1 g051(.A(KEYINPUT69), .B(new_n250_), .C1(new_n252_), .C2(new_n216_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n215_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n241_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n241_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n245_), .B1(new_n258_), .B2(KEYINPUT70), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n250_), .B1(new_n252_), .B2(new_n216_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n242_), .B1(new_n261_), .B2(new_n215_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n243_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n258_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G230gat), .A2(G233gat), .ZN(new_n265_));
  AND4_X1   g064(.A1(new_n246_), .A2(new_n260_), .A3(new_n264_), .A4(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(KEYINPUT67), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n241_), .B1(new_n233_), .B2(new_n243_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(new_n244_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n265_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n272_), .A2(KEYINPUT68), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT68), .B1(new_n272_), .B2(new_n273_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n267_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G120gat), .B(G148gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT5), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G176gat), .B(G204gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n272_), .A2(new_n273_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n272_), .A2(KEYINPUT68), .A3(new_n273_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n280_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n267_), .A3(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n281_), .A2(new_n288_), .A3(KEYINPUT71), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT71), .B1(new_n281_), .B2(new_n288_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT13), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n287_), .B1(new_n286_), .B2(new_n267_), .ZN(new_n294_));
  AOI211_X1 g093(.A(new_n266_), .B(new_n280_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n281_), .A2(new_n288_), .A3(KEYINPUT71), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT13), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n292_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT20), .ZN(new_n300_));
  INV_X1    g099(.A(G218gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G211gat), .ZN(new_n302_));
  INV_X1    g101(.A(G211gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G218gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT21), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G197gat), .A2(G204gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT92), .B(G204gat), .ZN(new_n309_));
  INV_X1    g108(.A(G197gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT93), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n306_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(KEYINPUT93), .B(new_n308_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT21), .ZN(new_n315_));
  INV_X1    g114(.A(G204gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT92), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT92), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G204gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n310_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n315_), .B1(new_n320_), .B2(new_n307_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(new_n319_), .A3(new_n310_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n315_), .B1(G197gat), .B2(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n305_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n313_), .A2(new_n314_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326_));
  INV_X1    g125(.A(G169gat), .ZN(new_n327_));
  INV_X1    g126(.A(G176gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT23), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G183gat), .A3(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n331_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT86), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n334_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n327_), .A2(new_n328_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(KEYINPUT24), .A3(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n335_), .A2(KEYINPUT86), .A3(G183gat), .A4(G190gat), .ZN(new_n344_));
  OR3_X1    g143(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n340_), .A2(new_n343_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT96), .ZN(new_n348_));
  INV_X1    g147(.A(G183gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT25), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G183gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n348_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n348_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT26), .B(G190gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n338_), .B1(new_n347_), .B2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n300_), .B1(new_n325_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n312_), .B1(new_n320_), .B2(new_n307_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n306_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n314_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n321_), .A2(new_n324_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n340_), .A2(new_n332_), .A3(new_n344_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n331_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n357_), .A2(new_n355_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n372_), .A2(new_n337_), .A3(new_n343_), .A4(new_n345_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n360_), .A2(new_n363_), .A3(new_n375_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n366_), .A2(new_n367_), .A3(new_n371_), .A4(new_n373_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT20), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT97), .B1(new_n325_), .B2(new_n359_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n337_), .A2(new_n332_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n370_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n350_), .A2(new_n352_), .A3(new_n348_), .ZN(new_n382_));
  XOR2_X1   g181(.A(KEYINPUT26), .B(G190gat), .Z(new_n383_));
  NOR3_X1   g182(.A1(new_n382_), .A2(new_n353_), .A3(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n381_), .B1(new_n384_), .B2(new_n346_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT97), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n368_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n378_), .B1(new_n379_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n376_), .B1(new_n388_), .B2(new_n363_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G8gat), .B(G36gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT18), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT98), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n393_), .B(new_n376_), .C1(new_n388_), .C2(new_n363_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n396_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n371_), .A2(new_n373_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n300_), .B1(new_n325_), .B2(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n368_), .A2(new_n386_), .A3(new_n385_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n386_), .B1(new_n368_), .B2(new_n385_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n362_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n393_), .B1(new_n405_), .B2(new_n376_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n399_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT27), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n398_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n388_), .A2(new_n363_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT20), .B1(new_n368_), .B2(new_n385_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n325_), .A2(new_n400_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n362_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(KEYINPUT27), .B(new_n397_), .C1(new_n414_), .C2(new_n393_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417_));
  INV_X1    g216(.A(G141gat), .ZN(new_n418_));
  INV_X1    g217(.A(G148gat), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .A4(KEYINPUT89), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT89), .ZN(new_n421_));
  OAI22_X1  g220(.A1(new_n421_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G141gat), .A2(G148gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT2), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n420_), .A2(new_n422_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(KEYINPUT1), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT1), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(G155gat), .A3(G162gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n434_), .A3(new_n428_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G141gat), .B(G148gat), .Z(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n431_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(KEYINPUT29), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G22gat), .B(G50gat), .Z(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n440_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n442_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT91), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(G228gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n447_), .A2(G228gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(G233gat), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n438_), .B2(KEYINPUT29), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n453_), .A2(new_n368_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n455_));
  NAND2_X1  g254(.A1(new_n438_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n451_), .B1(new_n368_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G78gat), .B(G106gat), .ZN(new_n458_));
  OR3_X1    g257(.A1(new_n454_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n458_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n460_));
  AND4_X1   g259(.A1(KEYINPUT95), .A2(new_n446_), .A3(new_n459_), .A4(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT95), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n463_), .A2(new_n446_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n416_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G71gat), .B(G99gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(G43gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n374_), .B(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G227gat), .A2(G233gat), .ZN(new_n471_));
  INV_X1    g270(.A(G15gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT30), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n470_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(KEYINPUT87), .ZN(new_n479_));
  XOR2_X1   g278(.A(G127gat), .B(G134gat), .Z(new_n480_));
  XOR2_X1   g279(.A(G113gat), .B(G120gat), .Z(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G127gat), .B(G134gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G113gat), .B(G120gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT31), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n478_), .A2(new_n479_), .A3(new_n487_), .ZN(new_n488_));
  OR3_X1    g287(.A1(new_n476_), .A2(new_n477_), .A3(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G57gat), .B(G85gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT103), .ZN(new_n492_));
  INV_X1    g291(.A(G1gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n495_));
  INV_X1    g294(.A(G29gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n494_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G225gat), .A2(G233gat), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n427_), .A2(new_n430_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n486_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT100), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n501_), .B2(new_n486_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n482_), .A2(new_n485_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n438_), .A2(new_n507_), .A3(new_n504_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT4), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT101), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n501_), .A2(new_n486_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NOR4_X1   g312(.A1(new_n501_), .A2(new_n486_), .A3(KEYINPUT101), .A4(KEYINPUT4), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n500_), .B1(new_n509_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n500_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n506_), .A2(new_n517_), .A3(new_n508_), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n499_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n499_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n490_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n467_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n399_), .A2(new_n406_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n411_), .A2(new_n412_), .A3(new_n362_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(new_n362_), .B2(new_n404_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n527_), .A2(new_n396_), .A3(new_n393_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT99), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT99), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n398_), .A2(new_n407_), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n509_), .A2(new_n500_), .A3(new_n515_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n517_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n532_), .A2(new_n498_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n520_), .A2(KEYINPUT33), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT33), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n499_), .B(new_n536_), .C1(new_n516_), .C2(new_n518_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n534_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n529_), .A2(new_n531_), .A3(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n393_), .A2(KEYINPUT32), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n410_), .A2(new_n413_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT104), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n527_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n527_), .B2(KEYINPUT104), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n521_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n465_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n416_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n465_), .A2(new_n521_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n490_), .B(KEYINPUT88), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n524_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G29gat), .B(G36gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT72), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G43gat), .B(G50gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n555_), .A2(KEYINPUT72), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(KEYINPUT72), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n559_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT79), .B(G15gat), .ZN(new_n569_));
  INV_X1    g368(.A(G22gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(G8gat), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT14), .B1(new_n493_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G1gat), .B(G8gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n568_), .A2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT84), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n563_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(KEYINPUT84), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .A4(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n576_), .B(new_n563_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(G229gat), .A3(G233gat), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(KEYINPUT85), .A3(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(KEYINPUT85), .B2(new_n582_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G169gat), .B(G197gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n586_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n299_), .A2(new_n554_), .A3(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G127gat), .B(G155gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT16), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT17), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n576_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n576_), .A2(new_n598_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n258_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n576_), .A2(new_n598_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n599_), .A3(new_n241_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n602_), .A2(KEYINPUT81), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT81), .B1(new_n602_), .B2(new_n604_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n597_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT82), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT82), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n609_), .B(new_n597_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n600_), .A2(new_n601_), .A3(new_n258_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n241_), .B1(new_n603_), .B2(new_n599_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n256_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n596_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n602_), .A2(KEYINPUT70), .A3(new_n604_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT80), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n614_), .A2(KEYINPUT80), .A3(new_n617_), .A4(new_n616_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n611_), .A2(KEYINPUT83), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT83), .B1(new_n611_), .B2(new_n622_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  OR2_X1    g424(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(KEYINPUT36), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n566_), .A2(new_n567_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n255_), .A2(KEYINPUT74), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT74), .ZN(new_n634_));
  INV_X1    g433(.A(new_n215_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n634_), .B1(new_n636_), .B2(new_n568_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  AOI22_X1  g437(.A1(new_n233_), .A2(new_n243_), .B1(new_n562_), .B2(new_n559_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT34), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(KEYINPUT35), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT75), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n563_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT75), .ZN(new_n645_));
  INV_X1    g444(.A(new_n642_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n638_), .A2(new_n643_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n641_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT35), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT76), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT74), .B1(new_n255_), .B2(new_n632_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n636_), .A2(new_n568_), .A3(new_n634_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n651_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n644_), .A2(new_n656_), .A3(new_n646_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n652_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n657_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n638_), .A3(KEYINPUT76), .ZN(new_n660_));
  AOI221_X4 g459(.A(new_n631_), .B1(new_n648_), .B2(new_n651_), .C1(new_n658_), .C2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n629_), .B(KEYINPUT36), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n658_), .A2(new_n660_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n648_), .A2(new_n651_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n626_), .B1(new_n661_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT78), .Z(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n626_), .B(new_n668_), .C1(new_n661_), .C2(new_n665_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n625_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n592_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n592_), .A2(KEYINPUT105), .A3(new_n673_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n521_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(G1gat), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT106), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n678_), .A2(new_n683_), .A3(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT38), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n550_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n466_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n553_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n523_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n661_), .A2(new_n665_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n611_), .A2(new_n622_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n299_), .A2(new_n591_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G1gat), .B1(new_n698_), .B2(new_n679_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n682_), .A2(KEYINPUT38), .A3(new_n684_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n687_), .A2(new_n699_), .A3(new_n700_), .ZN(G1324gat));
  INV_X1    g500(.A(KEYINPUT39), .ZN(new_n702_));
  INV_X1    g501(.A(new_n698_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(KEYINPUT107), .A3(new_n416_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(new_n698_), .B2(new_n548_), .ZN(new_n706_));
  AND4_X1   g505(.A1(new_n702_), .A2(new_n704_), .A3(G8gat), .A4(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n698_), .A2(new_n548_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n572_), .B1(new_n708_), .B2(KEYINPUT107), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n702_), .B1(new_n709_), .B2(new_n706_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n678_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n416_), .A2(new_n572_), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n707_), .A2(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT40), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI221_X1 g514(.A(KEYINPUT40), .B1(new_n711_), .B2(new_n712_), .C1(new_n707_), .C2(new_n710_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1325gat));
  NAND3_X1  g516(.A1(new_n678_), .A2(new_n472_), .A3(new_n552_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n719_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G15gat), .B1(new_n698_), .B2(new_n553_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT41), .Z(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n721_), .A3(new_n723_), .ZN(G1326gat));
  NAND3_X1  g523(.A1(new_n678_), .A2(new_n570_), .A3(new_n466_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G22gat), .B1(new_n698_), .B2(new_n465_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT42), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1327gat));
  NOR2_X1   g527(.A1(new_n623_), .A2(new_n624_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n693_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n592_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G29gat), .B1(new_n732_), .B2(new_n521_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n552_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n734_), .B(new_n672_), .C1(new_n735_), .C2(new_n524_), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n690_), .A2(new_n523_), .B1(new_n671_), .B2(new_n670_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n736_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n291_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n296_), .A2(KEYINPUT13), .A3(new_n297_), .ZN(new_n742_));
  AOI211_X1 g541(.A(new_n591_), .B(new_n729_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n740_), .A2(KEYINPUT44), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT111), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n625_), .B(new_n590_), .C1(new_n292_), .C2(new_n298_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n670_), .A2(new_n671_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n738_), .B1(new_n554_), .B2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n748_), .B2(new_n736_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(KEYINPUT44), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n745_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n740_), .A2(new_n743_), .ZN(new_n753_));
  XOR2_X1   g552(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n752_), .A2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n679_), .A2(new_n496_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n733_), .B1(new_n756_), .B2(new_n757_), .ZN(G1328gat));
  INV_X1    g557(.A(G36gat), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n592_), .A2(new_n759_), .A3(new_n416_), .A4(new_n730_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT45), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n548_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n762_));
  AOI211_X1 g561(.A(KEYINPUT112), .B(new_n759_), .C1(new_n752_), .C2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n750_), .B1(new_n749_), .B2(KEYINPUT44), .ZN(new_n765_));
  AND4_X1   g564(.A1(new_n750_), .A2(new_n740_), .A3(KEYINPUT44), .A4(new_n743_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n764_), .B1(new_n767_), .B2(G36gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n761_), .B1(new_n763_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT46), .B(new_n761_), .C1(new_n763_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1329gat));
  INV_X1    g572(.A(G43gat), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n490_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n752_), .A2(new_n755_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT113), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n752_), .A2(new_n778_), .A3(new_n755_), .A4(new_n775_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n774_), .B1(new_n731_), .B2(new_n553_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT47), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n777_), .A2(new_n783_), .A3(new_n779_), .A4(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1330gat));
  AOI21_X1  g584(.A(G50gat), .B1(new_n732_), .B2(new_n466_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n466_), .A2(G50gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n756_), .B2(new_n787_), .ZN(G1331gat));
  NAND2_X1  g587(.A1(new_n741_), .A2(new_n742_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n789_), .A2(new_n554_), .A3(new_n590_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n673_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(G57gat), .B1(new_n792_), .B2(new_n521_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT114), .ZN(new_n794_));
  NOR4_X1   g593(.A1(new_n694_), .A2(new_n789_), .A3(new_n625_), .A4(new_n590_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(G57gat), .A3(new_n521_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n794_), .A2(KEYINPUT115), .A3(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1332gat));
  INV_X1    g600(.A(G64gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n795_), .B2(new_n416_), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(KEYINPUT48), .Z(new_n804_));
  NAND3_X1  g603(.A1(new_n792_), .A2(new_n802_), .A3(new_n416_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1333gat));
  INV_X1    g605(.A(G71gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n795_), .B2(new_n552_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT116), .B(KEYINPUT49), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n792_), .A2(new_n807_), .A3(new_n552_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1334gat));
  NAND2_X1  g611(.A1(new_n795_), .A2(new_n466_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(G78gat), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n465_), .A2(G78gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n791_), .B2(new_n817_), .ZN(G1335gat));
  AND2_X1   g617(.A1(new_n790_), .A2(new_n730_), .ZN(new_n819_));
  AOI21_X1  g618(.A(G85gat), .B1(new_n819_), .B2(new_n521_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n789_), .A2(new_n729_), .A3(new_n590_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n740_), .A2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n822_), .A2(KEYINPUT118), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n822_), .A2(KEYINPUT118), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n521_), .A2(G85gat), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT119), .Z(new_n828_));
  AOI21_X1  g627(.A(new_n820_), .B1(new_n826_), .B2(new_n828_), .ZN(G1336gat));
  OAI21_X1  g628(.A(G92gat), .B1(new_n825_), .B2(new_n548_), .ZN(new_n830_));
  INV_X1    g629(.A(G92gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n819_), .A2(new_n831_), .A3(new_n416_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1337gat));
  OAI21_X1  g632(.A(G99gat), .B1(new_n825_), .B2(new_n553_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n490_), .A2(new_n208_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT120), .B1(new_n819_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT121), .B(KEYINPUT51), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1338gat));
  NAND3_X1  g638(.A1(new_n819_), .A2(new_n203_), .A3(new_n466_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n841_));
  INV_X1    g640(.A(new_n822_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n466_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n843_), .B2(G106gat), .ZN(new_n844_));
  AOI211_X1 g643(.A(KEYINPUT52), .B(new_n203_), .C1(new_n842_), .C2(new_n466_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n840_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n586_), .A2(new_n589_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n589_), .B1(new_n583_), .B2(new_n579_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n578_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n579_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n849_), .A2(new_n288_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n267_), .B2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n266_), .A2(KEYINPUT122), .A3(KEYINPUT55), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n267_), .A2(new_n855_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n268_), .A2(new_n271_), .A3(new_n246_), .A4(new_n260_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n273_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .A4(new_n860_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n861_), .A2(KEYINPUT56), .A3(new_n280_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT56), .B1(new_n861_), .B2(new_n280_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n853_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n747_), .B1(new_n848_), .B2(new_n864_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n864_), .A2(new_n848_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n590_), .B(new_n288_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n296_), .A2(new_n849_), .A3(new_n297_), .A4(new_n852_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n692_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT57), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n870_), .A2(KEYINPUT57), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n625_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n673_), .A2(new_n591_), .A3(new_n789_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT54), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  NOR4_X1   g677(.A1(new_n416_), .A2(new_n466_), .A3(new_n679_), .A4(new_n490_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n879_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n873_), .A2(KEYINPUT123), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n870_), .B2(KEYINPUT57), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n882_), .A2(new_n871_), .A3(new_n867_), .A4(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n695_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n881_), .B1(new_n886_), .B2(new_n876_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n880_), .B1(new_n887_), .B2(new_n878_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G113gat), .B1(new_n888_), .B2(new_n591_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n876_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n879_), .ZN(new_n891_));
  OR3_X1    g690(.A1(new_n891_), .A2(G113gat), .A3(new_n591_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n892_), .ZN(G1340gat));
  OAI21_X1  g692(.A(G120gat), .B1(new_n888_), .B2(new_n789_), .ZN(new_n894_));
  INV_X1    g693(.A(G120gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n789_), .B2(KEYINPUT60), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n887_), .B(new_n896_), .C1(KEYINPUT60), .C2(new_n895_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n897_), .ZN(G1341gat));
  OAI21_X1  g697(.A(G127gat), .B1(new_n888_), .B2(new_n695_), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n891_), .A2(G127gat), .A3(new_n625_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1342gat));
  OAI21_X1  g700(.A(G134gat), .B1(new_n888_), .B2(new_n747_), .ZN(new_n902_));
  OR3_X1    g701(.A1(new_n891_), .A2(G134gat), .A3(new_n693_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1343gat));
  NOR4_X1   g703(.A1(new_n552_), .A2(new_n679_), .A3(new_n465_), .A4(new_n416_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n890_), .A2(new_n590_), .A3(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g706(.A1(new_n890_), .A2(new_n299_), .A3(new_n905_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g708(.A1(new_n890_), .A2(new_n729_), .A3(new_n905_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT61), .B(G155gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1346gat));
  NAND2_X1  g711(.A1(new_n890_), .A2(new_n905_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G162gat), .B1(new_n913_), .B2(new_n747_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n693_), .A2(G162gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n913_), .B2(new_n915_), .ZN(G1347gat));
  NOR3_X1   g715(.A1(new_n553_), .A2(new_n521_), .A3(new_n466_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n416_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n919_), .A2(new_n326_), .A3(new_n590_), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n920_), .A2(KEYINPUT62), .A3(new_n327_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(KEYINPUT62), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n919_), .A2(new_n590_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n327_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n921_), .B1(new_n922_), .B2(new_n925_), .ZN(G1348gat));
  AOI21_X1  g725(.A(G176gat), .B1(new_n919_), .B2(new_n299_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n918_), .A2(new_n789_), .A3(new_n328_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n890_), .B2(new_n928_), .ZN(G1349gat));
  INV_X1    g728(.A(new_n918_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n729_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n886_), .B2(new_n876_), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n932_), .A2(KEYINPUT124), .ZN(new_n933_));
  AOI21_X1  g732(.A(G183gat), .B1(new_n932_), .B2(KEYINPUT124), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n695_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n933_), .A2(new_n934_), .B1(new_n919_), .B2(new_n935_), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n919_), .A2(new_n692_), .A3(new_n357_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n919_), .A2(new_n672_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n938_), .A2(new_n939_), .A3(G190gat), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(new_n938_), .B2(G190gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n937_), .B1(new_n940_), .B2(new_n941_), .ZN(G1351gat));
  NOR3_X1   g741(.A1(new_n552_), .A2(new_n521_), .A3(new_n465_), .ZN(new_n943_));
  OR2_X1    g742(.A1(new_n943_), .A2(KEYINPUT126), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(KEYINPUT126), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n944_), .A2(new_n416_), .A3(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n890_), .A2(new_n947_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949_), .B2(new_n590_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n948_), .A2(new_n310_), .A3(new_n591_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1352gat));
  NOR3_X1   g751(.A1(new_n948_), .A2(new_n309_), .A3(new_n789_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n949_), .A2(new_n299_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n953_), .B1(new_n316_), .B2(new_n954_), .ZN(G1353gat));
  NOR2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(KEYINPUT127), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n695_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n957_), .B1(new_n949_), .B2(new_n958_), .ZN(new_n959_));
  AND4_X1   g758(.A1(new_n890_), .A2(new_n947_), .A3(new_n957_), .A4(new_n958_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n959_), .A2(new_n960_), .ZN(G1354gat));
  OAI21_X1  g760(.A(G218gat), .B1(new_n948_), .B2(new_n747_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n692_), .A2(new_n301_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n962_), .B1(new_n948_), .B2(new_n963_), .ZN(G1355gat));
endmodule


