//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT21), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n202_), .A3(KEYINPUT21), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT22), .B(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(KEYINPUT81), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT23), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT79), .B(G190gat), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT78), .B(G183gat), .Z(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n215_), .A2(KEYINPUT81), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n216_), .A2(new_n217_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(KEYINPUT25), .ZN(new_n225_));
  OR2_X1    g024(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(KEYINPUT26), .ZN(new_n227_));
  OR2_X1    g026(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n228_));
  AOI22_X1  g027(.A1(new_n225_), .A2(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G169gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n213_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(KEYINPUT24), .A3(new_n217_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT80), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n231_), .A2(KEYINPUT80), .A3(KEYINPUT24), .A4(new_n217_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n219_), .A4(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n229_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n211_), .A2(new_n224_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT20), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n219_), .B1(G183gat), .B2(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n217_), .A2(KEYINPUT86), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n217_), .A2(KEYINPUT86), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n241_), .A2(new_n214_), .A3(new_n242_), .A4(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT25), .B(G183gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT26), .B(G190gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n247_), .A2(new_n219_), .A3(new_n236_), .A4(new_n232_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n240_), .B1(new_n249_), .B2(new_n210_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n239_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT19), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT85), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G8gat), .B(G36gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT18), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G64gat), .B(G92gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n211_), .B1(new_n238_), .B2(new_n224_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n253_), .ZN(new_n262_));
  OAI211_X1 g061(.A(KEYINPUT20), .B(new_n262_), .C1(new_n249_), .C2(new_n210_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n255_), .B(new_n260_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n251_), .A2(new_n254_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT20), .B1(new_n249_), .B2(new_n210_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT92), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT92), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n268_), .B(KEYINPUT20), .C1(new_n249_), .C2(new_n210_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n224_), .A2(new_n238_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n210_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n265_), .B1(new_n253_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n264_), .B1(new_n273_), .B2(new_n260_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT27), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT87), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n264_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n261_), .A2(new_n263_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n254_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n239_), .B2(new_n250_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n278_), .A2(new_n280_), .A3(new_n259_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT87), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n259_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n277_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n275_), .B1(KEYINPUT27), .B2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G155gat), .B(G162gat), .Z(new_n286_));
  OR3_X1    g085(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT83), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n287_), .B(new_n288_), .C1(new_n290_), .C2(KEYINPUT2), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n290_), .A2(KEYINPUT2), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n286_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n286_), .A2(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n295_), .A2(new_n289_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT84), .B(KEYINPUT29), .Z(new_n300_));
  OAI21_X1  g099(.A(new_n210_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(G228gat), .A3(G233gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G228gat), .A2(G233gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n303_), .B(new_n210_), .C1(new_n299_), .C2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G78gat), .B(G106gat), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n306_), .B(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n299_), .A2(new_n304_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G22gat), .B(G50gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n312_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n309_), .B(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n293_), .A2(new_n298_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G127gat), .B(G134gat), .Z(new_n318_));
  XOR2_X1   g117(.A(G113gat), .B(G120gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n317_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(KEYINPUT4), .ZN(new_n325_));
  INV_X1    g124(.A(new_n320_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n317_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n328_), .A2(KEYINPUT89), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(KEYINPUT89), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n324_), .B1(new_n331_), .B2(new_n323_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G1gat), .B(G29gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(G57gat), .B(G85gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n335_), .B(new_n336_), .Z(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n338_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n321_), .A2(KEYINPUT4), .B1(KEYINPUT89), .B2(new_n328_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n322_), .B1(new_n340_), .B2(new_n329_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n337_), .B1(new_n341_), .B2(new_n324_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G227gat), .A2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(G71gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(G99gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n270_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(new_n326_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G15gat), .B(G43gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT82), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT30), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT31), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n350_), .B(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n285_), .A2(new_n316_), .A3(new_n344_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT88), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n283_), .B1(new_n281_), .B2(KEYINPUT87), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n264_), .A2(new_n276_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT33), .B1(new_n332_), .B2(new_n338_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT33), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n362_), .B(new_n337_), .C1(new_n341_), .C2(new_n324_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT91), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n331_), .B2(new_n323_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n340_), .A2(KEYINPUT91), .A3(new_n322_), .A4(new_n329_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n337_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n277_), .A2(new_n282_), .A3(KEYINPUT88), .A4(new_n283_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n360_), .A2(new_n364_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT93), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n260_), .A2(KEYINPUT32), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n372_), .B1(new_n273_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n272_), .A2(new_n253_), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT93), .B(new_n375_), .C1(new_n376_), .C2(new_n265_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n255_), .B(new_n373_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n343_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n371_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n316_), .A2(new_n343_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n381_), .A2(new_n316_), .B1(new_n382_), .B2(new_n285_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n356_), .B1(new_n383_), .B2(new_n355_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G43gat), .B(G50gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G36gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G29gat), .ZN(new_n388_));
  INV_X1    g187(.A(G29gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G36gat), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n388_), .A2(new_n390_), .A3(KEYINPUT68), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT68), .B1(new_n388_), .B2(new_n390_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n386_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n390_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT68), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n388_), .A2(new_n390_), .A3(KEYINPUT68), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n385_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n393_), .A2(new_n398_), .A3(KEYINPUT15), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G15gat), .B(G22gat), .ZN(new_n400_));
  INV_X1    g199(.A(G1gat), .ZN(new_n401_));
  INV_X1    g200(.A(G8gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT14), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G8gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT73), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n405_), .A2(KEYINPUT73), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n404_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n405_), .A2(KEYINPUT73), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n410_), .A2(new_n403_), .A3(new_n400_), .A4(new_n406_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT15), .B1(new_n393_), .B2(new_n398_), .ZN(new_n413_));
  OR3_X1    g212(.A1(new_n399_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n393_), .A2(new_n398_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G229gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT76), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT75), .ZN(new_n420_));
  INV_X1    g219(.A(new_n415_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(new_n411_), .A3(new_n409_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n416_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n417_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n420_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  AOI211_X1 g224(.A(KEYINPUT75), .B(new_n417_), .C1(new_n422_), .C2(new_n416_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n419_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G113gat), .B(G141gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT77), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G169gat), .B(G197gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n419_), .B(new_n431_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n384_), .A2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n436_), .A2(KEYINPUT94), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(KEYINPUT94), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G85gat), .B(G92gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G99gat), .A2(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT6), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G99gat), .A3(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n440_), .B1(new_n444_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(G85gat), .B2(G92gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT9), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT65), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT65), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(new_n457_), .A3(new_n454_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n452_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT10), .B(G99gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n449_), .B1(new_n460_), .B2(G106gat), .ZN(new_n461_));
  OAI22_X1  g260(.A1(new_n450_), .A2(KEYINPUT8), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n440_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n466_));
  INV_X1    g265(.A(G99gat), .ZN(new_n467_));
  INV_X1    g266(.A(G106gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n441_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n470_), .A2(KEYINPUT66), .B1(new_n446_), .B2(new_n448_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT66), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n469_), .A2(new_n472_), .A3(new_n441_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n465_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  OAI22_X1  g273(.A1(new_n399_), .A2(new_n413_), .B1(new_n462_), .B2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n476_));
  NAND2_X1  g275(.A1(G232gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT35), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n470_), .A2(KEYINPUT66), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(new_n473_), .A3(new_n449_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n464_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n440_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n446_), .A2(new_n448_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(new_n470_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n463_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n456_), .A2(new_n458_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n452_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT10), .B(G99gat), .Z(new_n491_));
  AOI22_X1  g290(.A1(new_n491_), .A2(new_n468_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n421_), .A2(new_n483_), .A3(new_n487_), .A4(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n475_), .A2(new_n480_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT69), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT69), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n475_), .A2(new_n494_), .A3(new_n497_), .A4(new_n480_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G190gat), .B(G218gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G134gat), .B(G162gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n502_), .A2(KEYINPUT36), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n475_), .A2(new_n494_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n478_), .B(KEYINPUT35), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n499_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n496_), .A2(new_n498_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n502_), .B(KEYINPUT36), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n507_), .B(new_n508_), .C1(new_n509_), .C2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT71), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n499_), .A2(new_n506_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n515_), .A2(new_n516_), .A3(new_n508_), .A4(new_n507_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n510_), .B(KEYINPUT70), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n513_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n508_), .B1(new_n520_), .B2(new_n507_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT72), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n518_), .A2(new_n525_), .A3(new_n522_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT13), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT5), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT64), .Z(new_n535_));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G71gat), .B(G78gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT11), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(KEYINPUT11), .B2(new_n536_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n539_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(new_n462_), .B2(new_n474_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n545_));
  INV_X1    g344(.A(new_n537_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n538_), .B1(new_n547_), .B2(new_n541_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n483_), .A2(new_n548_), .A3(new_n487_), .A4(new_n493_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n544_), .A2(KEYINPUT12), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n551_), .B(new_n543_), .C1(new_n462_), .C2(new_n474_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n535_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n535_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n533_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n553_), .A2(new_n555_), .A3(new_n533_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n529_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n558_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(KEYINPUT13), .A3(new_n556_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G127gat), .B(G155gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT16), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G183gat), .B(G211gat), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  OR3_X1    g367(.A1(new_n567_), .A2(new_n568_), .A3(KEYINPUT17), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT17), .B1(new_n567_), .B2(new_n568_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT74), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n409_), .A2(new_n411_), .A3(new_n573_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n548_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n543_), .B1(new_n578_), .B2(new_n574_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n571_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n570_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n577_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n528_), .A2(new_n563_), .A3(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n439_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n401_), .A3(new_n343_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT38), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n356_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n381_), .A2(new_n316_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n382_), .A2(new_n285_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n355_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n590_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n515_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n507_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n435_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n563_), .A2(new_n600_), .A3(new_n584_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G1gat), .B1(new_n602_), .B2(new_n344_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n587_), .A2(new_n588_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n589_), .A2(new_n603_), .A3(new_n604_), .ZN(G1324gat));
  INV_X1    g404(.A(new_n285_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n586_), .A2(new_n402_), .A3(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G8gat), .B1(new_n602_), .B2(new_n285_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(KEYINPUT39), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(KEYINPUT39), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n607_), .B(KEYINPUT40), .C1(new_n610_), .C2(new_n609_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1325gat));
  OAI21_X1  g414(.A(G15gat), .B1(new_n602_), .B2(new_n594_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT95), .B(KEYINPUT41), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n616_), .A2(new_n617_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n586_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n594_), .A2(G15gat), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n618_), .B(new_n619_), .C1(new_n620_), .C2(new_n621_), .ZN(G1326gat));
  OAI21_X1  g421(.A(G22gat), .B1(new_n602_), .B2(new_n316_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT96), .Z(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(KEYINPUT42), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n620_), .A2(G22gat), .A3(new_n316_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(KEYINPUT42), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(G1327gat));
  INV_X1    g427(.A(new_n598_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n563_), .A2(new_n629_), .A3(new_n583_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n439_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n389_), .A3(new_n343_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n356_), .B(new_n634_), .C1(new_n383_), .C2(new_n355_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(KEYINPUT98), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n528_), .B(new_n635_), .C1(new_n595_), .C2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n384_), .A2(new_n528_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n636_), .A2(KEYINPUT97), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n636_), .A2(KEYINPUT97), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n638_), .A2(new_n641_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n563_), .A2(new_n600_), .A3(new_n583_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(KEYINPUT44), .A4(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n642_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n638_), .A3(new_n646_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT99), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n344_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G29gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n653_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n633_), .B1(new_n656_), .B2(new_n657_), .ZN(G1328gat));
  INV_X1    g457(.A(KEYINPUT46), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n285_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n387_), .B1(new_n652_), .B2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n285_), .A2(KEYINPUT101), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n285_), .A2(KEYINPUT101), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(G36gat), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n630_), .B(new_n666_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT45), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n659_), .B1(new_n661_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n649_), .A2(new_n650_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n606_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n651_), .B2(new_n647_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT46), .B(new_n668_), .C1(new_n673_), .C2(new_n387_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n674_), .ZN(G1329gat));
  NAND3_X1  g474(.A1(new_n671_), .A2(G43gat), .A3(new_n355_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n651_), .B2(new_n647_), .ZN(new_n677_));
  INV_X1    g476(.A(G43gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n678_), .B1(new_n631_), .B2(new_n594_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT47), .B1(new_n677_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT47), .ZN(new_n682_));
  INV_X1    g481(.A(new_n652_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n682_), .B(new_n679_), .C1(new_n683_), .C2(new_n676_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1330gat));
  OR3_X1    g484(.A1(new_n631_), .A2(G50gat), .A3(new_n316_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n316_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n652_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n687_), .B1(new_n652_), .B2(new_n688_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n686_), .B1(new_n690_), .B2(new_n691_), .ZN(G1331gat));
  NOR2_X1   g491(.A1(new_n562_), .A2(new_n435_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n384_), .A2(new_n583_), .A3(new_n629_), .A4(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n695_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G57gat), .B1(new_n699_), .B2(new_n344_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n384_), .A2(new_n693_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n583_), .A3(new_n527_), .ZN(new_n702_));
  OR3_X1    g501(.A1(new_n702_), .A2(G57gat), .A3(new_n344_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(G1332gat));
  OR3_X1    g503(.A1(new_n702_), .A2(G64gat), .A3(new_n665_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G64gat), .B1(new_n699_), .B2(new_n665_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT48), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT48), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(G1333gat));
  OAI21_X1  g508(.A(G71gat), .B1(new_n699_), .B2(new_n594_), .ZN(new_n710_));
  XOR2_X1   g509(.A(KEYINPUT104), .B(KEYINPUT49), .Z(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n710_), .A2(new_n712_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n355_), .A2(new_n346_), .ZN(new_n715_));
  OAI22_X1  g514(.A1(new_n713_), .A2(new_n714_), .B1(new_n702_), .B2(new_n715_), .ZN(G1334gat));
  OR3_X1    g515(.A1(new_n702_), .A2(G78gat), .A3(new_n316_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n316_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n696_), .A2(new_n697_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(G78gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G78gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n717_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1335gat));
  NOR3_X1   g524(.A1(new_n562_), .A2(new_n435_), .A3(new_n583_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n644_), .A2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G85gat), .B1(new_n727_), .B2(new_n344_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n701_), .A2(new_n584_), .A3(new_n598_), .ZN(new_n729_));
  INV_X1    g528(.A(G85gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n343_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n731_), .ZN(G1336gat));
  OAI21_X1  g531(.A(G92gat), .B1(new_n727_), .B2(new_n665_), .ZN(new_n733_));
  INV_X1    g532(.A(G92gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n729_), .A2(new_n734_), .A3(new_n606_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1337gat));
  OAI21_X1  g535(.A(G99gat), .B1(new_n727_), .B2(new_n594_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n729_), .A2(new_n355_), .A3(new_n491_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  XOR2_X1   g538(.A(KEYINPUT106), .B(KEYINPUT51), .Z(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(G1338gat));
  XNOR2_X1  g540(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n648_), .A2(new_n718_), .A3(new_n638_), .A4(new_n726_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n468_), .B1(new_n744_), .B2(KEYINPUT52), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT107), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n746_), .B(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n729_), .A2(new_n468_), .A3(new_n718_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n742_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n746_), .A2(new_n748_), .ZN(new_n752_));
  AOI22_X1  g551(.A1(new_n743_), .A2(new_n745_), .B1(KEYINPUT107), .B2(new_n747_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n750_), .B(new_n742_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n751_), .A2(new_n755_), .ZN(G1339gat));
  NOR2_X1   g555(.A1(new_n606_), .A2(new_n718_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n594_), .A2(new_n344_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n525_), .B1(new_n518_), .B2(new_n522_), .ZN(new_n761_));
  AOI211_X1 g560(.A(KEYINPUT72), .B(new_n521_), .C1(new_n512_), .C2(new_n517_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT58), .ZN(new_n763_));
  INV_X1    g562(.A(new_n418_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n414_), .A2(new_n416_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n431_), .B1(new_n423_), .B2(new_n418_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n434_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(new_n558_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n550_), .A2(new_n552_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n554_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n553_), .A2(KEYINPUT55), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT111), .B1(new_n771_), .B2(new_n554_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n550_), .A2(new_n552_), .A3(new_n777_), .A4(new_n535_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n774_), .A2(new_n775_), .A3(new_n776_), .A4(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n533_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n533_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n770_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n763_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n533_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n533_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n769_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(KEYINPUT113), .A3(KEYINPUT58), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n761_), .B(new_n762_), .C1(new_n786_), .C2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n558_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n434_), .B(new_n767_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n598_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT57), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT112), .B(KEYINPUT57), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n760_), .B1(new_n791_), .B2(new_n798_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n784_), .A2(new_n785_), .A3(new_n763_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT58), .B1(new_n789_), .B2(KEYINPUT113), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n524_), .B(new_n526_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n795_), .A2(new_n797_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n802_), .A2(KEYINPUT114), .A3(new_n796_), .A4(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n584_), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n433_), .A2(new_n583_), .A3(new_n434_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT109), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n433_), .A2(new_n583_), .A3(KEYINPUT109), .A4(new_n434_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(new_n559_), .A3(new_n561_), .A4(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n562_), .A2(KEYINPUT110), .A3(new_n808_), .A4(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n814_), .B(new_n815_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n527_), .B2(new_n814_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n759_), .B1(new_n805_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(G113gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n435_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n759_), .A2(KEYINPUT59), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n802_), .A2(new_n796_), .A3(new_n803_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n584_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n819_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(KEYINPUT116), .A3(new_n584_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n825_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT115), .B1(new_n821_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n583_), .B1(new_n826_), .B2(new_n760_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n819_), .B1(new_n835_), .B2(new_n804_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n834_), .B(KEYINPUT59), .C1(new_n836_), .C2(new_n759_), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n600_), .B(new_n831_), .C1(new_n833_), .C2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n823_), .B1(new_n838_), .B2(new_n822_), .ZN(G1340gat));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n562_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n821_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n562_), .B(new_n831_), .C1(new_n833_), .C2(new_n837_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n840_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n821_), .B2(new_n583_), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT117), .Z(new_n846_));
  NAND2_X1  g645(.A1(new_n833_), .A2(new_n837_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n831_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n847_), .A2(G127gat), .A3(new_n583_), .A4(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n846_), .A2(new_n849_), .ZN(G1342gat));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n527_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n831_), .B(new_n854_), .C1(new_n833_), .C2(new_n837_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G134gat), .B1(new_n821_), .B2(new_n598_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n851_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n847_), .A2(new_n848_), .A3(new_n853_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n856_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(KEYINPUT118), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n857_), .A2(new_n860_), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n836_), .A2(new_n355_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n664_), .A2(new_n316_), .A3(new_n344_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n805_), .A2(new_n820_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n594_), .A3(new_n864_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT119), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n600_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT120), .B(G141gat), .Z(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1344gat));
  AOI21_X1  g670(.A(new_n562_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT121), .B(G148gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1345gat));
  AOI21_X1  g673(.A(new_n584_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n875_), .B(new_n877_), .ZN(G1346gat));
  NAND2_X1  g677(.A1(new_n865_), .A2(new_n868_), .ZN(new_n879_));
  INV_X1    g678(.A(G162gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(new_n598_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n527_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n880_), .ZN(G1347gat));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n829_), .A2(new_n830_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n355_), .A2(new_n344_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n665_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n718_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n885_), .A2(new_n435_), .A3(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n885_), .A2(new_n212_), .A3(new_n435_), .A4(new_n889_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT62), .B1(new_n890_), .B2(G169gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n884_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n894_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n896_), .A2(KEYINPUT122), .A3(new_n892_), .A4(new_n891_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1348gat));
  NAND3_X1  g697(.A1(new_n885_), .A2(new_n563_), .A3(new_n889_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n836_), .A2(new_n718_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n888_), .A2(new_n213_), .A3(new_n562_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n899_), .A2(new_n213_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT123), .Z(G1349gat));
  NAND3_X1  g702(.A1(new_n900_), .A2(new_n583_), .A3(new_n887_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n221_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n885_), .A2(new_n889_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n584_), .A2(new_n245_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n904_), .A2(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(G1350gat));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n528_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G190gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n906_), .A2(new_n246_), .A3(new_n598_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1351gat));
  XOR2_X1   g711(.A(KEYINPUT124), .B(G197gat), .Z(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n664_), .A2(new_n382_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n862_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n600_), .ZN(new_n917_));
  MUX2_X1   g716(.A(new_n913_), .B(new_n914_), .S(new_n917_), .Z(G1352gat));
  INV_X1    g717(.A(new_n916_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n562_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922_));
  INV_X1    g721(.A(G204gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(KEYINPUT125), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n921_), .B(new_n924_), .ZN(G1353gat));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  AND2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n916_), .A2(new_n584_), .A3(new_n926_), .A4(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n919_), .A2(new_n583_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n926_), .ZN(G1354gat));
  AND3_X1   g729(.A1(new_n919_), .A2(G218gat), .A3(new_n528_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n916_), .A2(new_n629_), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n932_), .A2(KEYINPUT127), .ZN(new_n933_));
  AOI21_X1  g732(.A(G218gat), .B1(new_n932_), .B2(KEYINPUT127), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n931_), .B1(new_n933_), .B2(new_n934_), .ZN(G1355gat));
endmodule


