//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(G113gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(G120gat), .Z(new_n205_));
  XOR2_X1   g004(.A(new_n205_), .B(KEYINPUT31), .Z(new_n206_));
  NAND2_X1  g005(.A1(G227gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(G15gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G71gat), .B(G99gat), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n208_), .B(new_n209_), .Z(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT80), .ZN(new_n212_));
  AOI21_X1  g011(.A(G176gat), .B1(new_n212_), .B2(KEYINPUT22), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT81), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(G169gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT23), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(G183gat), .B2(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(G169gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT78), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT79), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n222_), .A2(KEYINPUT24), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n229_), .A2(new_n217_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n222_), .A2(new_n231_), .A3(KEYINPUT24), .A4(new_n223_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n225_), .A2(new_n226_), .A3(new_n230_), .A4(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT30), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n220_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n220_), .B2(new_n233_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n236_), .A2(G43gat), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G43gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n220_), .A2(new_n233_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT30), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n241_), .B2(new_n235_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n211_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(G43gat), .B1(new_n236_), .B2(new_n237_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n239_), .A3(new_n235_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n210_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT82), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT82), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n243_), .A2(new_n249_), .A3(new_n246_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n206_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT83), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n252_), .B1(new_n247_), .B2(new_n206_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  AOI211_X1 g053(.A(new_n252_), .B(new_n206_), .C1(new_n248_), .C2(new_n250_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT27), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(G36gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G64gat), .B(G92gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT92), .B(G8gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n228_), .B(KEYINPUT88), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n227_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT24), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n221_), .A2(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n266_), .A2(new_n217_), .A3(new_n224_), .A4(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT22), .B(G169gat), .ZN(new_n270_));
  INV_X1    g069(.A(G176gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n218_), .A2(new_n223_), .A3(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n273_), .A2(KEYINPUT89), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(KEYINPUT89), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n269_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G197gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G204gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT86), .B(G204gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT21), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G211gat), .B(G218gat), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G197gat), .A2(G204gat), .ZN(new_n284_));
  OAI211_X1 g083(.A(KEYINPUT21), .B(new_n284_), .C1(new_n279_), .C2(G197gat), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n285_), .B(new_n282_), .C1(new_n280_), .C2(KEYINPUT21), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n276_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n287_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(new_n220_), .A3(new_n233_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(KEYINPUT20), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT19), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT90), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT90), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(new_n296_), .A3(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n276_), .A2(new_n287_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n293_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n240_), .A2(new_n287_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n299_), .A2(KEYINPUT20), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n264_), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n291_), .A2(new_n296_), .A3(new_n293_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n296_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n264_), .B(new_n302_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n257_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n289_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n309_), .A2(new_n301_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n300_), .B1(new_n310_), .B2(KEYINPUT20), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n291_), .A2(new_n293_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n263_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n306_), .A2(KEYINPUT27), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  INV_X1    g117(.A(G155gat), .ZN(new_n319_));
  INV_X1    g118(.A(G162gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n319_), .A2(new_n320_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n324_), .B(KEYINPUT84), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n323_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT85), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n317_), .B(new_n318_), .C1(new_n325_), .C2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n322_), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n316_), .B(KEYINPUT3), .Z(new_n330_));
  XOR2_X1   g129(.A(new_n318_), .B(KEYINPUT2), .Z(new_n331_));
  OAI211_X1 g130(.A(new_n329_), .B(new_n321_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT29), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n287_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n335_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n339_), .B2(new_n289_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G78gat), .B(G106gat), .Z(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n336_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n333_), .A2(KEYINPUT29), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G22gat), .B(G50gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT28), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n347_), .B(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n342_), .B1(new_n336_), .B2(new_n340_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n346_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G1gat), .B(G29gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G57gat), .B(G85gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n205_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n333_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT93), .B1(new_n363_), .B2(KEYINPUT4), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n328_), .A2(new_n205_), .A3(new_n332_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(KEYINPUT4), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT93), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n333_), .A2(new_n369_), .A3(new_n362_), .A4(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n364_), .A2(new_n366_), .A3(new_n368_), .A4(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n363_), .A2(new_n367_), .A3(new_n365_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n361_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n373_), .A3(new_n361_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NOR4_X1   g176(.A1(new_n256_), .A2(new_n315_), .A3(new_n355_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n298_), .A2(new_n379_), .A3(new_n302_), .ZN(new_n380_));
  OAI211_X1 g179(.A(KEYINPUT32), .B(new_n264_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n376_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n380_), .B(new_n381_), .C1(new_n382_), .C2(new_n374_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n302_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n263_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .A4(new_n371_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n363_), .A2(new_n368_), .A3(new_n365_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n360_), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n306_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT33), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n376_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n372_), .A2(KEYINPUT33), .A3(new_n373_), .A4(new_n361_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n354_), .B(new_n383_), .C1(new_n389_), .C2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT27), .B1(new_n385_), .B2(new_n306_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n306_), .A2(new_n313_), .A3(KEYINPUT27), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n377_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n394_), .B(new_n256_), .C1(new_n397_), .C2(new_n354_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT95), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n248_), .A2(new_n250_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n206_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(KEYINPUT83), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(new_n253_), .B2(new_n251_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n377_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n308_), .A2(new_n404_), .A3(new_n314_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n405_), .B2(new_n355_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT95), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n394_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n378_), .B1(new_n399_), .B2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT74), .B(G1gat), .Z(new_n410_));
  INV_X1    g209(.A(G8gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT14), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G15gat), .B(G22gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(G1gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G8gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT69), .B(G29gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G36gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(G43gat), .B(G50gat), .Z(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n415_), .B(new_n411_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n418_), .A2(new_n419_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n418_), .A2(new_n419_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G229gat), .A2(G233gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n421_), .A2(new_n426_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n429_), .B1(new_n428_), .B2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G113gat), .B(G141gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G169gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(new_n277_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n428_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n438_), .B1(new_n442_), .B2(new_n429_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G230gat), .A2(G233gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AND3_X1   g246(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT9), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G85gat), .B(G92gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(G99gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT10), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT10), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G99gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(G106gat), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G92gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n451_), .A2(KEYINPUT64), .A3(G85gat), .ZN(new_n460_));
  OR2_X1    g259(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n453_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT65), .ZN(new_n464_));
  INV_X1    g263(.A(G106gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n454_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT7), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT7), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n464_), .A2(new_n468_), .A3(new_n454_), .A4(new_n465_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n450_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n452_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT8), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT8), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n463_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G57gat), .ZN(new_n477_));
  INV_X1    g276(.A(G64gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G57gat), .A2(G64gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G71gat), .B(G78gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT11), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n479_), .A2(new_n485_), .A3(new_n480_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n481_), .A2(new_n483_), .A3(KEYINPUT11), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT66), .B1(new_n476_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n459_), .A2(G85gat), .ZN(new_n491_));
  INV_X1    g290(.A(G85gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G92gat), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n451_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n462_), .A2(new_n494_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n458_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n470_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n474_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n502_), .B(new_n489_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT66), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n490_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n476_), .A2(new_n489_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n447_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n512_));
  NOR4_X1   g311(.A1(new_n453_), .A2(KEYINPUT67), .A3(new_n458_), .A4(new_n462_), .ZN(new_n513_));
  OAI22_X1  g312(.A1(new_n512_), .A2(new_n513_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n489_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(KEYINPUT12), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT12), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n476_), .B2(new_n489_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n516_), .A2(new_n518_), .A3(new_n446_), .A4(new_n505_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n510_), .A2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G120gat), .B(G148gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G204gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT5), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G176gat), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n520_), .A2(new_n524_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(new_n528_), .B2(KEYINPUT13), .ZN(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n530_));
  NAND3_X1  g329(.A1(new_n525_), .A2(new_n526_), .A3(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n445_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n409_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G190gat), .B(G218gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(G134gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n320_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT36), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT71), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n420_), .A2(new_n431_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n433_), .A2(new_n542_), .A3(new_n514_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT34), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n476_), .A2(new_n420_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n546_), .A2(new_n547_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n541_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n552_), .A2(new_n539_), .A3(new_n538_), .A4(new_n553_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT73), .B1(new_n557_), .B2(KEYINPUT37), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n554_), .A2(KEYINPUT72), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n556_), .B1(new_n554_), .B2(KEYINPUT72), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT37), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  OAI211_X1 g361(.A(KEYINPUT73), .B(KEYINPUT37), .C1(new_n559_), .C2(new_n560_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G127gat), .B(G155gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT76), .ZN(new_n567_));
  XOR2_X1   g366(.A(G183gat), .B(G211gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n489_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n416_), .B(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n571_), .B1(new_n574_), .B2(KEYINPUT77), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT17), .Z(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n571_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n565_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n535_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n377_), .A3(new_n410_), .ZN(new_n582_));
  XOR2_X1   g381(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n557_), .B(KEYINPUT97), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n578_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n535_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G1gat), .B1(new_n589_), .B2(new_n404_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n590_), .ZN(G1324gat));
  AOI21_X1  g390(.A(new_n411_), .B1(new_n588_), .B2(new_n315_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT39), .Z(new_n593_));
  NAND3_X1  g392(.A1(new_n581_), .A2(new_n411_), .A3(new_n315_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT40), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(G1325gat));
  INV_X1    g396(.A(G15gat), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n588_), .B2(new_n403_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT41), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n581_), .A2(new_n598_), .A3(new_n403_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1326gat));
  INV_X1    g401(.A(G22gat), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n588_), .B2(new_n355_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT42), .Z(new_n605_));
  NAND3_X1  g404(.A1(new_n581_), .A2(new_n603_), .A3(new_n355_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(G1327gat));
  INV_X1    g406(.A(new_n578_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(new_n585_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n535_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT101), .ZN(new_n611_));
  INV_X1    g410(.A(G29gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n377_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n564_), .B(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT43), .B1(new_n409_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n378_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n398_), .A2(KEYINPUT95), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n407_), .B1(new_n406_), .B2(new_n394_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n564_), .A2(KEYINPUT43), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AOI211_X1 g421(.A(new_n608_), .B(new_n534_), .C1(new_n616_), .C2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT100), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n608_), .B1(new_n616_), .B2(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n533_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(KEYINPUT44), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT100), .B(new_n631_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n404_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n613_), .B1(new_n633_), .B2(new_n612_), .ZN(G1328gat));
  INV_X1    g433(.A(KEYINPUT46), .ZN(new_n635_));
  INV_X1    g434(.A(G36gat), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n629_), .A2(KEYINPUT44), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n628_), .B1(new_n627_), .B2(KEYINPUT99), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n632_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n636_), .B1(new_n639_), .B2(new_n315_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n611_), .A2(new_n636_), .A3(new_n315_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT45), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n635_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n641_), .B(KEYINPUT45), .ZN(new_n645_));
  INV_X1    g444(.A(new_n315_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n645_), .B(KEYINPUT46), .C1(new_n636_), .C2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(G1329gat));
  AOI211_X1 g448(.A(new_n239_), .B(new_n256_), .C1(new_n630_), .C2(new_n632_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n611_), .A2(new_n403_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(KEYINPUT102), .A2(G43gat), .ZN(new_n652_));
  OR2_X1    g451(.A1(KEYINPUT102), .A2(G43gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT47), .B1(new_n650_), .B2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n639_), .A2(G43gat), .A3(new_n403_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT47), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n654_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(new_n659_), .ZN(G1330gat));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n661_));
  INV_X1    g460(.A(G50gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n639_), .B2(new_n355_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n611_), .A2(new_n662_), .A3(new_n355_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n354_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT103), .B(new_n664_), .C1(new_n667_), .C2(new_n662_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1331gat));
  NAND2_X1  g468(.A1(new_n620_), .A2(new_n445_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(new_n532_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n579_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n477_), .B1(new_n674_), .B2(new_n404_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT105), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT105), .ZN(new_n677_));
  INV_X1    g476(.A(new_n532_), .ZN(new_n678_));
  NOR4_X1   g477(.A1(new_n670_), .A2(new_n586_), .A3(new_n578_), .A4(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(G57gat), .A3(new_n377_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT106), .Z(new_n681_));
  NOR3_X1   g480(.A1(new_n676_), .A2(new_n677_), .A3(new_n681_), .ZN(G1332gat));
  AOI21_X1  g481(.A(new_n478_), .B1(new_n679_), .B2(new_n315_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT48), .Z(new_n684_));
  NAND2_X1  g483(.A1(new_n315_), .A2(new_n478_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n674_), .B2(new_n685_), .ZN(G1333gat));
  INV_X1    g485(.A(G71gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n679_), .B2(new_n403_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT49), .Z(new_n689_));
  NAND2_X1  g488(.A1(new_n403_), .A2(new_n687_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n674_), .B2(new_n690_), .ZN(G1334gat));
  INV_X1    g490(.A(G78gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n679_), .B2(new_n355_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT107), .B(KEYINPUT108), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT50), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n693_), .B(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n354_), .A2(G78gat), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT109), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n674_), .B2(new_n698_), .ZN(G1335gat));
  NAND3_X1  g498(.A1(new_n626_), .A2(new_n445_), .A3(new_n532_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n701_));
  AOI211_X1 g500(.A(new_n404_), .B(new_n700_), .C1(new_n461_), .C2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n673_), .A2(new_n609_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n492_), .B1(new_n703_), .B2(new_n404_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n704_), .A2(KEYINPUT110), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(KEYINPUT110), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1336gat));
  INV_X1    g506(.A(new_n703_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n459_), .A3(new_n315_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G92gat), .B1(new_n700_), .B2(new_n646_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT111), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n713_), .A3(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1337gat));
  INV_X1    g514(.A(new_n455_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n457_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n708_), .A2(new_n719_), .A3(new_n403_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G99gat), .B1(new_n700_), .B2(new_n256_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT51), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n720_), .A2(new_n724_), .A3(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1338gat));
  INV_X1    g525(.A(KEYINPUT53), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n626_), .A2(new_n355_), .A3(new_n445_), .A4(new_n532_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G106gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT52), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n729_), .A2(new_n732_), .A3(G106gat), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n354_), .A2(G106gat), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n672_), .A2(new_n532_), .A3(new_n609_), .A4(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n728_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n729_), .A2(new_n732_), .A3(G106gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n732_), .B1(new_n729_), .B2(G106gat), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n728_), .B(new_n736_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n727_), .B1(new_n737_), .B2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT112), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(KEYINPUT53), .A3(new_n740_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n742_), .A2(new_n745_), .ZN(G1339gat));
  NOR3_X1   g545(.A1(new_n578_), .A2(KEYINPUT113), .A3(new_n444_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(new_n532_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT113), .B1(new_n578_), .B2(new_n444_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n564_), .A3(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT54), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n516_), .B(new_n518_), .C1(new_n490_), .C2(new_n507_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n752_), .A2(KEYINPUT115), .A3(new_n447_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT115), .B1(new_n752_), .B2(new_n447_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n519_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT114), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n519_), .A2(new_n758_), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n753_), .A2(new_n754_), .B1(new_n756_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT116), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n519_), .A2(new_n755_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n519_), .B2(new_n758_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n763_), .B(new_n764_), .C1(new_n754_), .C2(new_n753_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n524_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n761_), .A2(KEYINPUT56), .A3(new_n524_), .A4(new_n765_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n761_), .A2(new_n765_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n772_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n524_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n771_), .A2(new_n444_), .A3(new_n525_), .A4(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT118), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n434_), .A2(new_n441_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n776_), .B(new_n438_), .C1(new_n441_), .C2(new_n427_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n440_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n527_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n766_), .A2(new_n769_), .A3(new_n767_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n525_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n444_), .A4(new_n771_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n775_), .A2(new_n779_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT57), .B1(new_n785_), .B2(new_n585_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT119), .B(KEYINPUT57), .C1(new_n785_), .C2(new_n585_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n785_), .A2(KEYINPUT57), .A3(new_n585_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n781_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n778_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n778_), .A2(new_n791_), .A3(KEYINPUT58), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n565_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n790_), .A2(new_n796_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n788_), .A2(new_n789_), .A3(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n751_), .B1(new_n798_), .B2(new_n608_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n646_), .A2(new_n377_), .A3(new_n354_), .A4(new_n403_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT120), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT59), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n578_), .B1(new_n797_), .B2(new_n786_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n751_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n801_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n803_), .A2(G113gat), .A3(new_n444_), .A4(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n203_), .B1(new_n802_), .B2(new_n445_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1340gat));
  XOR2_X1   g609(.A(KEYINPUT121), .B(G120gat), .Z(new_n811_));
  AND2_X1   g610(.A1(new_n532_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n799_), .B(new_n801_), .C1(KEYINPUT60), .C2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n803_), .A2(new_n813_), .A3(new_n532_), .A4(new_n807_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n811_), .B1(new_n813_), .B2(KEYINPUT60), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1341gat));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n817_));
  OAI21_X1  g616(.A(G127gat), .B1(new_n578_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(G127gat), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT122), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n803_), .A2(new_n807_), .A3(new_n818_), .A4(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n802_), .B2(new_n578_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1342gat));
  NAND4_X1  g622(.A1(new_n803_), .A2(G134gat), .A3(new_n565_), .A4(new_n807_), .ZN(new_n824_));
  INV_X1    g623(.A(G134gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n802_), .B2(new_n585_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1343gat));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n750_), .B(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n785_), .A2(new_n585_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT119), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n790_), .A2(new_n796_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n786_), .A2(new_n787_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n829_), .B1(new_n836_), .B2(new_n578_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n837_), .A2(new_n354_), .A3(new_n403_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n315_), .A2(new_n404_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OR3_X1    g639(.A1(new_n840_), .A2(G141gat), .A3(new_n445_), .ZN(new_n841_));
  OAI21_X1  g640(.A(G141gat), .B1(new_n840_), .B2(new_n445_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1344gat));
  AND2_X1   g642(.A1(new_n838_), .A2(new_n839_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT123), .B(G148gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n532_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n845_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n840_), .B2(new_n678_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1345gat));
  XNOR2_X1  g648(.A(KEYINPUT61), .B(G155gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n844_), .B2(new_n608_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n850_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n840_), .A2(new_n578_), .A3(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1346gat));
  AOI21_X1  g653(.A(G162gat), .B1(new_n844_), .B2(new_n586_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n840_), .A2(new_n320_), .A3(new_n615_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1347gat));
  XNOR2_X1  g656(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n646_), .A2(new_n377_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n256_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n355_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n805_), .A2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(G169gat), .B1(new_n865_), .B2(new_n445_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT125), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n868_), .B(G169gat), .C1(new_n865_), .C2(new_n445_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n859_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n858_), .B1(new_n866_), .B2(KEYINPUT125), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n444_), .A2(new_n270_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(KEYINPUT126), .Z(new_n873_));
  OAI22_X1  g672(.A1(new_n870_), .A2(new_n871_), .B1(new_n865_), .B2(new_n873_), .ZN(G1348gat));
  INV_X1    g673(.A(new_n865_), .ZN(new_n875_));
  AOI21_X1  g674(.A(G176gat), .B1(new_n875_), .B2(new_n532_), .ZN(new_n876_));
  NOR4_X1   g675(.A1(new_n837_), .A2(new_n271_), .A3(new_n355_), .A4(new_n863_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n532_), .ZN(G1349gat));
  NOR3_X1   g677(.A1(new_n865_), .A2(new_n578_), .A3(new_n227_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n799_), .A2(new_n608_), .A3(new_n354_), .A4(new_n862_), .ZN(new_n880_));
  INV_X1    g679(.A(G183gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(G1350gat));
  OAI21_X1  g681(.A(G190gat), .B1(new_n865_), .B2(new_n564_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n586_), .A2(new_n265_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n865_), .B2(new_n884_), .ZN(G1351gat));
  NAND4_X1  g684(.A1(new_n799_), .A2(new_n355_), .A3(new_n256_), .A4(new_n860_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n445_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n277_), .ZN(G1352gat));
  NOR4_X1   g687(.A1(new_n837_), .A2(new_n354_), .A3(new_n403_), .A4(new_n861_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n532_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G204gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n279_), .B2(new_n890_), .ZN(G1353gat));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n893_));
  INV_X1    g692(.A(G211gat), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n578_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n889_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n897_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n886_), .A2(KEYINPUT127), .A3(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n895_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n889_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT127), .B1(new_n886_), .B2(new_n899_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(new_n893_), .A4(new_n894_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(G1354gat));
  AND3_X1   g704(.A1(new_n889_), .A2(G218gat), .A3(new_n565_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G218gat), .B1(new_n889_), .B2(new_n586_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1355gat));
endmodule


