//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n563_,
    new_n564_, new_n565_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT37), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT68), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT15), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G92gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(KEYINPUT9), .A3(new_n215_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n217_), .A2(KEYINPUT67), .A3(new_n221_), .A4(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n214_), .A2(new_n221_), .A3(new_n225_), .A4(new_n216_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n215_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AOI211_X1 g035(.A(KEYINPUT8), .B(new_n232_), .C1(new_n236_), .C2(new_n214_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT8), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT7), .ZN(new_n239_));
  INV_X1    g038(.A(G99gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n219_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n212_), .B1(G99gat), .B2(G106gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n233_), .B(new_n241_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n232_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n238_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n237_), .A2(new_n246_), .A3(KEYINPUT66), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n211_), .A2(new_n213_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n241_), .A2(new_n233_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n245_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT8), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n244_), .A2(new_n238_), .A3(new_n245_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n248_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n231_), .B1(new_n247_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n209_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n227_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n208_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT35), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G190gat), .B(G218gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G134gat), .B(G162gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n260_), .A2(new_n261_), .B1(KEYINPUT36), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G232gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(new_n260_), .B2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n256_), .A2(KEYINPUT69), .A3(new_n259_), .A4(new_n268_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n264_), .A2(KEYINPUT36), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n265_), .A2(new_n271_), .A3(new_n276_), .A4(new_n272_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n203_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n277_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n278_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G15gat), .B(G22gat), .ZN(new_n284_));
  INV_X1    g083(.A(G1gat), .ZN(new_n285_));
  INV_X1    g084(.A(G8gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT14), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G1gat), .B(G8gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G231gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G57gat), .B(G64gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G71gat), .B(G78gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT11), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(KEYINPUT11), .ZN(new_n296_));
  INV_X1    g095(.A(new_n294_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n293_), .A2(KEYINPUT11), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n295_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n292_), .B(new_n300_), .Z(new_n301_));
  XNOR2_X1  g100(.A(G127gat), .B(G155gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT16), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G183gat), .B(G211gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT17), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT71), .Z(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT72), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n305_), .B(KEYINPUT17), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n301_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n283_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT73), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n209_), .A2(new_n290_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n290_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n208_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G229gat), .A2(G233gat), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n315_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n208_), .B(new_n316_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n318_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G113gat), .B(G141gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT74), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n324_), .B(KEYINPUT75), .Z(new_n325_));
  XNOR2_X1  g124(.A(G169gat), .B(G197gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  OR3_X1    g126(.A1(new_n319_), .A2(new_n322_), .A3(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n327_), .B1(new_n319_), .B2(new_n322_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT23), .ZN(new_n334_));
  INV_X1    g133(.A(G169gat), .ZN(new_n335_));
  INV_X1    g134(.A(G176gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n334_), .B1(KEYINPUT24), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT24), .B1(new_n335_), .B2(new_n336_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT77), .B(KEYINPUT25), .Z(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G183gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT78), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n345_), .A3(G183gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT26), .B(G190gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT76), .B(G183gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT25), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n344_), .A2(new_n346_), .A3(new_n347_), .A4(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n341_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n348_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n334_), .B1(new_n352_), .B2(G190gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(G169gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G197gat), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n358_), .A2(KEYINPUT83), .A3(G204gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(G197gat), .B(G204gat), .Z(new_n360_));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n361_));
  OAI211_X1 g160(.A(KEYINPUT21), .B(new_n359_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G211gat), .B(G218gat), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n362_), .B(new_n363_), .C1(KEYINPUT21), .C2(new_n360_), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(KEYINPUT84), .Z(new_n365_));
  INV_X1    g164(.A(KEYINPUT21), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n360_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n367_), .B2(new_n360_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n364_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n332_), .B1(new_n357_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n340_), .A2(KEYINPUT88), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT88), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n339_), .A2(new_n376_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n338_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT25), .B(G183gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT87), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n347_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT22), .B(G169gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT89), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n336_), .ZN(new_n385_));
  OR2_X1    g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n334_), .A2(new_n386_), .B1(G169gat), .B2(G176gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n382_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n371_), .B(new_n374_), .C1(new_n370_), .C2(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n357_), .A2(new_n370_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n332_), .B1(new_n389_), .B2(new_n370_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT90), .B1(new_n393_), .B2(new_n373_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT90), .ZN(new_n395_));
  AOI211_X1 g194(.A(new_n395_), .B(new_n374_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n390_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT18), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n401_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n403_), .B(new_n390_), .C1(new_n394_), .C2(new_n396_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT27), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n393_), .A2(new_n373_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n370_), .A2(KEYINPUT86), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n370_), .A2(KEYINPUT86), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n382_), .A4(new_n388_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n374_), .B1(new_n411_), .B2(new_n371_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n401_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n404_), .A2(KEYINPUT27), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n407_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G127gat), .B(G134gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT79), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G113gat), .B(G120gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n417_), .B(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G155gat), .B(G162gat), .Z(new_n421_));
  INV_X1    g220(.A(KEYINPUT1), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n424_));
  OR2_X1    g223(.A1(G141gat), .A2(G148gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G141gat), .A2(G148gat), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n428_), .B(KEYINPUT80), .Z(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(KEYINPUT81), .ZN(new_n430_));
  AOI22_X1  g229(.A1(KEYINPUT2), .A2(new_n430_), .B1(new_n425_), .B2(KEYINPUT3), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(KEYINPUT2), .B2(new_n430_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n421_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n420_), .A2(new_n427_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n427_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n417_), .B(new_n418_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT91), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n435_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(KEYINPUT91), .A3(new_n420_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT4), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n444_), .B(KEYINPUT92), .Z(new_n445_));
  OR2_X1    g244(.A1(new_n437_), .A2(KEYINPUT4), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n445_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n442_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G1gat), .B(G29gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G85gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT0), .B(G57gat), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n452_), .B(new_n453_), .Z(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n447_), .A2(new_n454_), .A3(new_n449_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G71gat), .B(G99gat), .ZN(new_n460_));
  INV_X1    g259(.A(G43gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n357_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(new_n420_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465_));
  INV_X1    g264(.A(G15gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT30), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT31), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n464_), .B(new_n469_), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n459_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT29), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n440_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT82), .B(KEYINPUT28), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G228gat), .A2(G233gat), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n477_), .B(new_n370_), .C1(new_n440_), .C2(new_n472_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n409_), .A2(new_n410_), .B1(KEYINPUT29), .B2(new_n435_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n477_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n475_), .B(new_n478_), .C1(new_n477_), .C2(new_n479_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G78gat), .B(G106gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(G22gat), .B(G50gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n481_), .A2(new_n482_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n415_), .A2(new_n471_), .A3(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n407_), .A2(new_n459_), .A3(new_n488_), .A4(new_n414_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n457_), .A2(KEYINPUT33), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n457_), .A2(KEYINPUT33), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n443_), .A2(new_n448_), .A3(new_n446_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n454_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n402_), .A2(new_n496_), .A3(new_n404_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n403_), .A2(KEYINPUT32), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT94), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n498_), .B(KEYINPUT93), .Z(new_n501_));
  OAI211_X1 g300(.A(new_n501_), .B(new_n390_), .C1(new_n394_), .C2(new_n396_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n503_), .B(new_n498_), .C1(new_n408_), .C2(new_n412_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n500_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n493_), .A2(new_n497_), .B1(new_n505_), .B2(new_n458_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n490_), .B1(new_n506_), .B2(new_n488_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n470_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n489_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G230gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT64), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n300_), .B(new_n227_), .C1(new_n237_), .C2(new_n246_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT65), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n258_), .A2(KEYINPUT65), .A3(new_n300_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n258_), .A2(new_n300_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n511_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n258_), .B2(new_n300_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n511_), .B1(new_n258_), .B2(new_n300_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT66), .B1(new_n237_), .B2(new_n246_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n252_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n230_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n300_), .A2(new_n519_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n520_), .B(new_n521_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n518_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G120gat), .B(G148gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT5), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G176gat), .B(G204gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n531_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n518_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(KEYINPUT13), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(KEYINPUT13), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NOR4_X1   g338(.A1(new_n314_), .A2(new_n331_), .A3(new_n509_), .A4(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT95), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(new_n285_), .A3(new_n458_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT38), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n543_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n509_), .A2(new_n280_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n539_), .A2(new_n331_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n312_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT96), .Z(new_n550_));
  AND2_X1   g349(.A1(new_n546_), .A2(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n551_), .A2(new_n458_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n544_), .B(new_n545_), .C1(new_n285_), .C2(new_n552_), .ZN(G1324gat));
  NAND3_X1  g352(.A1(new_n541_), .A2(new_n286_), .A3(new_n415_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n551_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n415_), .ZN(new_n556_));
  OAI21_X1  g355(.A(G8gat), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(KEYINPUT39), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(KEYINPUT39), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n554_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT40), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(G1325gat));
  NAND3_X1  g361(.A1(new_n541_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n466_), .B1(new_n551_), .B2(new_n470_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT41), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(G1326gat));
  INV_X1    g365(.A(G22gat), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n541_), .A2(new_n567_), .A3(new_n488_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n551_), .B2(new_n488_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT97), .B(KEYINPUT42), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(G1327gat));
  NOR2_X1   g371(.A1(new_n509_), .A2(new_n331_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n280_), .A2(new_n312_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(new_n539_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n576_), .A2(G29gat), .A3(new_n459_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT43), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n275_), .A2(new_n277_), .A3(new_n282_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n280_), .B2(new_n203_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n578_), .B1(new_n509_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n488_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n402_), .A2(new_n496_), .A3(new_n404_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n492_), .B2(new_n491_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n500_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n459_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n582_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n470_), .B1(new_n587_), .B2(new_n490_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT43), .B(new_n283_), .C1(new_n588_), .C2(new_n489_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n581_), .A2(new_n589_), .A3(new_n312_), .A4(new_n547_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT44), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n591_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n458_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n577_), .B1(new_n594_), .B2(G29gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT98), .Z(G1328gat));
  NOR2_X1   g395(.A1(new_n556_), .A2(G36gat), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n573_), .A2(new_n575_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(KEYINPUT99), .B(KEYINPUT45), .Z(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n599_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n592_), .A2(new_n415_), .A3(new_n593_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(G36gat), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(G1329gat));
  NAND4_X1  g409(.A1(new_n592_), .A2(G43gat), .A3(new_n470_), .A4(new_n593_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n461_), .B1(new_n576_), .B2(new_n508_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g413(.A1(new_n592_), .A2(G50gat), .A3(new_n488_), .A4(new_n593_), .ZN(new_n615_));
  INV_X1    g414(.A(G50gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n576_), .B2(new_n582_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n615_), .A2(new_n617_), .ZN(G1331gat));
  INV_X1    g417(.A(new_n539_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n548_), .A2(new_n331_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n546_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G57gat), .B1(new_n623_), .B2(new_n459_), .ZN(new_n624_));
  NOR4_X1   g423(.A1(new_n314_), .A2(new_n330_), .A3(new_n509_), .A4(new_n619_), .ZN(new_n625_));
  INV_X1    g424(.A(G57gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n458_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(G1332gat));
  NOR2_X1   g427(.A1(new_n556_), .A2(G64gat), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT104), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n625_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G64gat), .B1(new_n623_), .B2(new_n556_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT103), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT102), .B(KEYINPUT48), .Z(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n633_), .A2(new_n635_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n631_), .B1(new_n636_), .B2(new_n637_), .ZN(G1333gat));
  INV_X1    g437(.A(G71gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n622_), .B2(new_n470_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT49), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n625_), .A2(new_n639_), .A3(new_n470_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1334gat));
  INV_X1    g442(.A(G78gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n622_), .B2(new_n488_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n625_), .A2(new_n644_), .A3(new_n488_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1335gat));
  NOR4_X1   g448(.A1(new_n509_), .A2(new_n330_), .A3(new_n619_), .A4(new_n574_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(new_n222_), .A3(new_n458_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n283_), .B1(new_n588_), .B2(new_n489_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n548_), .B1(new_n652_), .B2(new_n578_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n619_), .A2(new_n330_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n653_), .A2(KEYINPUT106), .A3(new_n589_), .A4(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n581_), .A2(new_n589_), .A3(new_n312_), .A4(new_n654_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n459_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n651_), .B1(new_n659_), .B2(new_n222_), .ZN(G1336gat));
  NAND3_X1  g459(.A1(new_n650_), .A2(new_n223_), .A3(new_n415_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n556_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n661_), .B1(new_n662_), .B2(new_n223_), .ZN(G1337gat));
  NAND4_X1  g462(.A1(new_n650_), .A2(new_n470_), .A3(new_n218_), .A4(new_n220_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n655_), .A2(new_n658_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n470_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT107), .B1(new_n666_), .B2(G99gat), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n668_), .B(new_n240_), .C1(new_n665_), .C2(new_n470_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n664_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT51), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT51), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n672_), .B(new_n664_), .C1(new_n667_), .C2(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(G1338gat));
  NAND3_X1  g473(.A1(new_n650_), .A2(new_n219_), .A3(new_n488_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n656_), .A2(new_n582_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT52), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(G106gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(new_n676_), .B2(G106gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g481(.A1(new_n415_), .A2(new_n488_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n458_), .A3(new_n470_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT59), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n330_), .A2(new_n534_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n526_), .A2(KEYINPUT55), .ZN(new_n689_));
  INV_X1    g488(.A(new_n525_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n255_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT55), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n691_), .A2(new_n692_), .A3(new_n520_), .A4(new_n521_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n520_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n511_), .B1(new_n694_), .B2(new_n516_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT109), .B(new_n511_), .C1(new_n694_), .C2(new_n516_), .ZN(new_n698_));
  AOI221_X4 g497(.A(KEYINPUT110), .B1(new_n689_), .B2(new_n693_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n698_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n693_), .A2(new_n689_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n531_), .B1(new_n699_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT56), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n691_), .A2(new_n514_), .A3(new_n515_), .A4(new_n520_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT109), .B1(new_n707_), .B2(new_n511_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n698_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n702_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT110), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n701_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(KEYINPUT56), .A3(new_n531_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n688_), .B1(new_n706_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n320_), .A2(new_n318_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n327_), .A2(new_n716_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n717_), .A2(KEYINPUT111), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n315_), .A2(new_n317_), .A3(new_n321_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(KEYINPUT111), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n721_), .A2(new_n328_), .A3(new_n535_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n279_), .B1(new_n715_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT57), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n721_), .A2(new_n328_), .A3(new_n534_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT56), .B1(new_n713_), .B2(new_n531_), .ZN(new_n728_));
  AOI211_X1 g527(.A(new_n705_), .B(new_n533_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT58), .B(new_n727_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT58), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n580_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n730_), .A2(new_n733_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n726_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n723_), .A2(new_n724_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n731_), .A2(new_n732_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n730_), .A3(new_n283_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(KEYINPUT112), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n312_), .B1(new_n736_), .B2(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n620_), .A2(new_n539_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT108), .B(KEYINPUT54), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n580_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n743_), .B2(new_n580_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n687_), .B1(new_n742_), .B2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n312_), .B1(new_n740_), .B2(new_n725_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n749_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n686_), .B1(new_n752_), .B2(new_n685_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT113), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n734_), .A2(new_n726_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n748_), .B1(new_n755_), .B2(new_n312_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT59), .B1(new_n756_), .B2(new_n684_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n725_), .B1(new_n740_), .B2(KEYINPUT112), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n734_), .A2(new_n735_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n748_), .B1(new_n761_), .B2(new_n312_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n757_), .B(new_n758_), .C1(new_n762_), .C2(new_n687_), .ZN(new_n763_));
  INV_X1    g562(.A(G113gat), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n331_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n754_), .A2(new_n763_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n752_), .A2(new_n685_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n764_), .B1(new_n767_), .B2(new_n331_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n766_), .A2(KEYINPUT114), .A3(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1340gat));
  OAI21_X1  g572(.A(new_n757_), .B1(new_n762_), .B2(new_n687_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G120gat), .B1(new_n774_), .B2(new_n619_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT60), .ZN(new_n776_));
  AOI21_X1  g575(.A(G120gat), .B1(new_n539_), .B2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT115), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n776_), .B2(G120gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n752_), .A2(new_n685_), .A3(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT116), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n775_), .A2(new_n781_), .ZN(G1341gat));
  INV_X1    g581(.A(G127gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n767_), .B2(new_n312_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT117), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n754_), .A2(new_n763_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n312_), .A2(new_n783_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n786_), .B2(new_n787_), .ZN(G1342gat));
  NAND3_X1  g587(.A1(new_n754_), .A2(new_n763_), .A3(new_n283_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(G134gat), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n279_), .A2(G134gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n767_), .B2(new_n791_), .ZN(G1343gat));
  NOR2_X1   g591(.A1(new_n582_), .A2(new_n470_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n556_), .A2(new_n458_), .A3(new_n793_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT118), .Z(new_n795_));
  NAND2_X1  g594(.A1(new_n752_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n331_), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g597(.A1(new_n796_), .A2(new_n619_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT119), .B(G148gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(G1345gat));
  NOR2_X1   g600(.A1(new_n796_), .A2(new_n312_), .ZN(new_n802_));
  XOR2_X1   g601(.A(KEYINPUT61), .B(G155gat), .Z(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(G1346gat));
  OAI21_X1  g603(.A(G162gat), .B1(new_n796_), .B2(new_n580_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n279_), .A2(G162gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n796_), .B2(new_n806_), .ZN(G1347gat));
  NOR2_X1   g606(.A1(new_n556_), .A2(new_n471_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n488_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n548_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n330_), .B(new_n810_), .C1(new_n811_), .C2(new_n748_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G169gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n742_), .A2(new_n749_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(new_n330_), .A3(new_n384_), .A4(new_n810_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(KEYINPUT62), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT62), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n812_), .A2(new_n818_), .A3(G169gat), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n816_), .A2(new_n817_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n817_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1348gat));
  AND2_X1   g621(.A1(new_n814_), .A2(new_n810_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G176gat), .B1(new_n823_), .B2(new_n539_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n756_), .A2(new_n488_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n809_), .A2(new_n336_), .A3(new_n619_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(G1349gat));
  NOR2_X1   g626(.A1(new_n809_), .A2(new_n312_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n352_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n312_), .A2(new_n380_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n823_), .B2(new_n830_), .ZN(G1350gat));
  NAND2_X1  g630(.A1(new_n280_), .A2(new_n347_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT121), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n823_), .A2(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n823_), .A2(new_n283_), .ZN(new_n835_));
  INV_X1    g634(.A(G190gat), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT122), .B(new_n834_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838_));
  INV_X1    g637(.A(new_n834_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n836_), .B1(new_n823_), .B2(new_n283_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n841_), .ZN(G1351gat));
  NAND3_X1  g641(.A1(new_n793_), .A2(new_n459_), .A3(new_n415_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n752_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n358_), .B1(new_n845_), .B2(new_n331_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT124), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n848_), .B(new_n358_), .C1(new_n845_), .C2(new_n331_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n752_), .A2(G197gat), .A3(new_n330_), .A4(new_n844_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT123), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT125), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT125), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n850_), .A2(new_n855_), .A3(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1352gat));
  NOR2_X1   g656(.A1(new_n845_), .A2(new_n619_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT126), .B(G204gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1353gat));
  INV_X1    g659(.A(KEYINPUT63), .ZN(new_n861_));
  INV_X1    g660(.A(G211gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n548_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT127), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n752_), .A2(new_n844_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n861_), .A2(new_n862_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1354gat));
  OAI21_X1  g666(.A(G218gat), .B1(new_n845_), .B2(new_n580_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n279_), .A2(G218gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n845_), .B2(new_n869_), .ZN(G1355gat));
endmodule


