//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n829_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202_));
  AOI21_X1  g001(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206_));
  OAI22_X1  g005(.A1(new_n203_), .A2(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(new_n204_), .B2(new_n203_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n205_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(KEYINPUT3), .B2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT82), .Z(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n214_), .B(KEYINPUT1), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n209_), .B(new_n216_), .C1(new_n212_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G197gat), .B(G204gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G211gat), .B(G218gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT84), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n223_), .B(new_n226_), .Z(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT85), .B(KEYINPUT21), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT86), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n227_), .B1(new_n224_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G228gat), .A2(G233gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n220_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT87), .ZN(new_n235_));
  INV_X1    g034(.A(new_n219_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n232_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n233_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT87), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n220_), .A2(new_n241_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n235_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G78gat), .B(G106gat), .Z(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n202_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT28), .B(G22gat), .ZN(new_n248_));
  INV_X1    g047(.A(G50gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n247_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT90), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT90), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n246_), .A2(new_n254_), .A3(new_n251_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n243_), .B(new_n244_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n253_), .A2(new_n257_), .A3(new_n255_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G225gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT78), .ZN(new_n265_));
  INV_X1    g064(.A(G113gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G120gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT79), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n267_), .B(G120gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT79), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(new_n273_), .A3(new_n219_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n269_), .A2(new_n236_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n275_), .B1(new_n274_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n263_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n278_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(new_n263_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G1gat), .B(G29gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G85gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT0), .ZN(new_n287_));
  INV_X1    g086(.A(G57gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n280_), .A2(new_n283_), .A3(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT25), .B(G183gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n298_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n296_), .A2(KEYINPUT76), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT76), .B1(new_n296_), .B2(new_n299_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT23), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(KEYINPUT24), .B2(new_n297_), .ZN(new_n304_));
  OR3_X1    g103(.A1(new_n300_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(G183gat), .B2(G190gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G169gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n232_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n304_), .B(KEYINPUT91), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n296_), .A2(new_n299_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n309_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n311_), .B(KEYINPUT20), .C1(new_n232_), .C2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT19), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n232_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n320_), .B(KEYINPUT20), .C1(new_n232_), .C2(new_n310_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G8gat), .B(G36gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT18), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G64gat), .ZN(new_n325_));
  INV_X1    g124(.A(G92gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT32), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n322_), .A2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n315_), .A2(new_n317_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n321_), .A2(new_n317_), .ZN(new_n331_));
  OAI211_X1 g130(.A(KEYINPUT32), .B(new_n327_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n293_), .A2(new_n329_), .A3(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n262_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n334_), .B(new_n290_), .C1(new_n262_), .C2(new_n281_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT93), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n292_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n322_), .A2(new_n327_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n327_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n319_), .B(new_n340_), .C1(new_n318_), .C2(new_n321_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(KEYINPUT92), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT92), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n322_), .A2(new_n343_), .A3(new_n327_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n280_), .A2(new_n283_), .A3(KEYINPUT33), .A4(new_n289_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n338_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n261_), .B(new_n333_), .C1(new_n336_), .C2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350_));
  INV_X1    g149(.A(G43gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT30), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G227gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n310_), .B(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT77), .B(G15gat), .Z(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n356_), .A2(new_n357_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n354_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n310_), .B(new_n355_), .Z(new_n362_));
  INV_X1    g161(.A(new_n357_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(new_n353_), .A3(new_n358_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(KEYINPUT80), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT31), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT31), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n361_), .A2(KEYINPUT80), .A3(new_n368_), .A4(new_n365_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n270_), .A2(new_n273_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n367_), .A2(new_n270_), .A3(new_n273_), .A4(new_n369_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n372_), .A2(KEYINPUT81), .A3(new_n373_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n340_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n339_), .A2(KEYINPUT27), .A3(new_n378_), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n379_), .A2(KEYINPUT94), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(KEYINPUT94), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n342_), .A2(new_n382_), .A3(new_n344_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(new_n293_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n376_), .B(new_n377_), .C1(new_n261_), .C2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT95), .B1(new_n349_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n376_), .A2(new_n377_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT95), .ZN(new_n390_));
  INV_X1    g189(.A(new_n261_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n293_), .B2(new_n384_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n389_), .A2(new_n390_), .A3(new_n348_), .A4(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n293_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT96), .B1(new_n391_), .B2(new_n384_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n384_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT96), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n261_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n374_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n387_), .A2(new_n393_), .B1(new_n394_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G230gat), .A2(G233gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n401_), .B(KEYINPUT64), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT9), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(KEYINPUT66), .ZN(new_n405_));
  INV_X1    g204(.A(G85gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n326_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G85gat), .A2(G92gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT9), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n404_), .A2(KEYINPUT66), .ZN(new_n412_));
  AND2_X1   g211(.A1(G85gat), .A2(G92gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G99gat), .A2(G106gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT6), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(G99gat), .A3(G106gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT65), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT10), .B(G99gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(G106gat), .ZN(new_n423_));
  INV_X1    g222(.A(G106gat), .ZN(new_n424_));
  INV_X1    g223(.A(G99gat), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n425_), .A2(KEYINPUT10), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(KEYINPUT10), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT65), .B(new_n424_), .C1(new_n426_), .C2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n415_), .A2(new_n420_), .A3(new_n423_), .A4(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n407_), .A2(new_n408_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n417_), .A2(new_n419_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT7), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(new_n425_), .A3(new_n424_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n430_), .B1(new_n431_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT8), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n420_), .A2(new_n434_), .A3(new_n433_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(KEYINPUT8), .A3(new_n430_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n429_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G57gat), .B(G64gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G71gat), .B(G78gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n446_));
  XOR2_X1   g245(.A(G71gat), .B(G78gat), .Z(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(KEYINPUT11), .A3(new_n442_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n445_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n441_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n449_), .A2(new_n429_), .A3(new_n438_), .A4(new_n440_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(KEYINPUT12), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT12), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n441_), .A2(new_n454_), .A3(new_n450_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n403_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n451_), .A2(new_n458_), .A3(new_n452_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n441_), .A2(KEYINPUT67), .A3(new_n450_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n403_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n457_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G120gat), .B(G148gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT5), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(G176gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G204gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n462_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT13), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT15), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(G43gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n249_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n472_), .B(new_n351_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(G50gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n471_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(G50gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n249_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(KEYINPUT15), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G1gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT71), .B(G22gat), .ZN(new_n483_));
  INV_X1    g282(.A(G15gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT72), .B(G1gat), .Z(new_n486_));
  INV_X1    g285(.A(G8gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n482_), .B1(new_n485_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(new_n482_), .A3(new_n488_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(G8gat), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n491_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n487_), .B1(new_n493_), .B2(new_n489_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n481_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n478_), .A2(new_n479_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n496_), .B1(new_n494_), .B2(new_n492_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT75), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n481_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT75), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n497_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n494_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(KEYINPUT74), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n499_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT74), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n494_), .A2(new_n508_), .A3(new_n496_), .A4(new_n492_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n506_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G113gat), .B(G141gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(G169gat), .ZN(new_n512_));
  INV_X1    g311(.A(G197gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n503_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n503_), .B2(new_n510_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n470_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n400_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n441_), .A2(new_n496_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n481_), .B2(new_n441_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT34), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT35), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n526_), .A2(new_n527_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n523_), .A2(new_n527_), .A3(new_n526_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT68), .B(KEYINPUT36), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G190gat), .B(G218gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G134gat), .ZN(new_n536_));
  INV_X1    g335(.A(G162gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(KEYINPUT36), .Z(new_n540_));
  OAI21_X1  g339(.A(new_n539_), .B1(new_n533_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT37), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n529_), .A2(new_n530_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n532_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(KEYINPUT69), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n533_), .A2(KEYINPUT69), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n539_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n542_), .B(KEYINPUT70), .C1(KEYINPUT37), .C2(new_n549_), .ZN(new_n550_));
  OR3_X1    g349(.A1(new_n549_), .A2(KEYINPUT70), .A3(KEYINPUT37), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n494_), .A2(new_n492_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n449_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n553_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G127gat), .B(G155gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT16), .ZN(new_n560_));
  INV_X1    g359(.A(G183gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(G211gat), .ZN(new_n563_));
  OR3_X1    g362(.A1(new_n557_), .A2(new_n558_), .A3(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(KEYINPUT17), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n557_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT73), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n552_), .A2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n521_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n293_), .A3(new_n486_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT38), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n571_), .B1(KEYINPUT98), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(KEYINPUT98), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n387_), .A2(new_n393_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n399_), .A2(new_n394_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n519_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n549_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n579_), .A2(new_n580_), .A3(new_n567_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n581_), .A2(KEYINPUT97), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(KEYINPUT97), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n293_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(G1gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n575_), .A2(new_n585_), .ZN(G1324gat));
  NAND3_X1  g385(.A1(new_n581_), .A2(KEYINPUT100), .A3(new_n384_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n567_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n521_), .A2(new_n549_), .A3(new_n384_), .A4(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT100), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n587_), .A2(G8gat), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT39), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n587_), .A2(KEYINPUT39), .A3(G8gat), .A4(new_n591_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n570_), .A2(new_n487_), .A3(new_n384_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT99), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n570_), .A2(new_n598_), .A3(new_n487_), .A4(new_n384_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n594_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT40), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n594_), .A2(new_n600_), .A3(KEYINPUT40), .A4(new_n595_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(G1325gat));
  NAND3_X1  g404(.A1(new_n570_), .A2(new_n484_), .A3(new_n388_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n582_), .A2(new_n388_), .A3(new_n583_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n607_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT41), .B1(new_n607_), .B2(G15gat), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n606_), .B1(new_n608_), .B2(new_n609_), .ZN(G1326gat));
  INV_X1    g409(.A(G22gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n261_), .B(KEYINPUT101), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n570_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n582_), .A2(new_n583_), .A3(new_n612_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT42), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n614_), .A2(new_n615_), .A3(G22gat), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n614_), .B2(G22gat), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n613_), .B1(new_n616_), .B2(new_n617_), .ZN(G1327gat));
  NAND3_X1  g417(.A1(new_n578_), .A2(KEYINPUT43), .A3(new_n552_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT43), .ZN(new_n620_));
  INV_X1    g419(.A(new_n552_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n620_), .B1(new_n400_), .B2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n619_), .A2(new_n622_), .A3(new_n519_), .A4(new_n568_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT44), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n624_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n293_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT102), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n623_), .B(KEYINPUT44), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n293_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n631_), .A3(G29gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n568_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n549_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT103), .Z(new_n635_));
  NOR2_X1   g434(.A1(new_n579_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n293_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n638_), .ZN(G1328gat));
  INV_X1    g438(.A(KEYINPUT46), .ZN(new_n640_));
  INV_X1    g439(.A(G36gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n629_), .B2(new_n384_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n636_), .A2(new_n641_), .A3(new_n384_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT45), .Z(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n625_), .A2(new_n384_), .A3(new_n626_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G36gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n643_), .B(KEYINPUT45), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(KEYINPUT46), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n645_), .A2(new_n649_), .ZN(G1329gat));
  NOR2_X1   g449(.A1(new_n374_), .A2(new_n351_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n629_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n636_), .A2(new_n388_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n351_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT47), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT47), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n652_), .A2(new_n657_), .A3(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1330gat));
  NAND3_X1  g458(.A1(new_n625_), .A2(new_n391_), .A3(new_n626_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT104), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n629_), .A2(new_n662_), .A3(new_n391_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n663_), .A3(G50gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n636_), .A2(new_n249_), .A3(new_n612_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1331gat));
  INV_X1    g465(.A(new_n518_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n400_), .A2(new_n667_), .A3(new_n469_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(new_n569_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G57gat), .B1(new_n669_), .B2(new_n293_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n549_), .A3(new_n633_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n671_), .A2(new_n288_), .A3(new_n394_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1332gat));
  NOR2_X1   g472(.A1(new_n396_), .A2(G64gat), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT105), .Z(new_n675_));
  NAND2_X1  g474(.A1(new_n669_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G64gat), .B1(new_n671_), .B2(new_n396_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT48), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT48), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT106), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n676_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1333gat));
  OAI21_X1  g483(.A(G71gat), .B1(new_n671_), .B2(new_n389_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT49), .ZN(new_n686_));
  INV_X1    g485(.A(G71gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n669_), .A2(new_n687_), .A3(new_n388_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1334gat));
  NAND4_X1  g488(.A1(new_n668_), .A2(new_n549_), .A3(new_n633_), .A4(new_n612_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G78gat), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT50), .ZN(new_n692_));
  INV_X1    g491(.A(G78gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n669_), .A2(new_n693_), .A3(new_n612_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1335gat));
  INV_X1    g494(.A(new_n635_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n668_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n293_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n469_), .A2(new_n667_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n619_), .A2(new_n622_), .A3(new_n568_), .A4(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n394_), .A2(new_n406_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n698_), .B1(new_n702_), .B2(new_n703_), .ZN(G1336gat));
  AOI21_X1  g503(.A(G92gat), .B1(new_n697_), .B2(new_n384_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n396_), .A2(new_n326_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n702_), .B2(new_n706_), .ZN(G1337gat));
  AOI21_X1  g506(.A(new_n425_), .B1(new_n702_), .B2(new_n388_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n374_), .A2(new_n422_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n697_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT108), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT51), .B1(new_n708_), .B2(new_n711_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n700_), .A2(KEYINPUT107), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n700_), .A2(KEYINPUT107), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n388_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G99gat), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n716_), .A2(KEYINPUT108), .A3(new_n717_), .A4(new_n710_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n712_), .A2(new_n718_), .ZN(G1338gat));
  NAND4_X1  g518(.A1(new_n668_), .A2(new_n424_), .A3(new_n391_), .A4(new_n696_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT109), .Z(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT52), .B(G106gat), .C1(new_n700_), .C2(new_n261_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G106gat), .B1(new_n700_), .B2(new_n261_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n721_), .A2(new_n722_), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT53), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT53), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n721_), .A2(new_n728_), .A3(new_n725_), .A4(new_n722_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1339gat));
  NAND2_X1  g529(.A1(new_n453_), .A2(new_n455_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT112), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n453_), .A2(new_n733_), .A3(new_n455_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n403_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT113), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT114), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n456_), .B2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT55), .B1(new_n456_), .B2(new_n737_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n732_), .A2(new_n742_), .A3(new_n403_), .A4(new_n734_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n737_), .B(KEYINPUT55), .C1(new_n456_), .C2(new_n738_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n736_), .A2(new_n741_), .A3(new_n743_), .A4(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n467_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(KEYINPUT56), .A3(new_n467_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n462_), .A2(new_n467_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n498_), .A2(new_n507_), .A3(new_n502_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n506_), .A2(new_n499_), .A3(new_n509_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n514_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT115), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n503_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n753_), .A2(new_n754_), .A3(new_n758_), .A4(new_n514_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n756_), .A2(new_n757_), .A3(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n750_), .A2(new_n752_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT58), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n750_), .A2(KEYINPUT58), .A3(new_n752_), .A4(new_n760_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n552_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766_));
  INV_X1    g565(.A(new_n517_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n751_), .B1(new_n767_), .B2(new_n757_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n749_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT56), .B1(new_n745_), .B2(new_n467_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n760_), .A2(new_n468_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n580_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n766_), .B(KEYINPUT57), .C1(new_n773_), .C2(KEYINPUT116), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n752_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n776_));
  AND4_X1   g575(.A1(new_n757_), .A2(new_n756_), .A3(new_n468_), .A4(new_n759_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n549_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT117), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n778_), .B2(KEYINPUT117), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n765_), .B(new_n774_), .C1(new_n780_), .C2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT118), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n567_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n552_), .A2(new_n667_), .A3(new_n568_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n469_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n786_), .A2(new_n469_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT54), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n786_), .A2(KEYINPUT110), .A3(new_n787_), .A4(new_n469_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n785_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n399_), .A2(new_n293_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G113gat), .B1(new_n799_), .B2(new_n667_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n783_), .A2(new_n568_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n783_), .A2(KEYINPUT119), .A3(new_n568_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n794_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n798_), .A2(KEYINPUT59), .B1(new_n807_), .B2(new_n797_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n518_), .A2(new_n266_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n800_), .B1(new_n808_), .B2(new_n809_), .ZN(G1340gat));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n470_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT60), .B1(new_n470_), .B2(new_n268_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n798_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(G120gat), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n798_), .A2(new_n812_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(KEYINPUT60), .B2(new_n815_), .ZN(G1341gat));
  AOI21_X1  g615(.A(G127gat), .B1(new_n799_), .B2(new_n633_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n588_), .A2(G127gat), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT120), .Z(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n808_), .B2(new_n819_), .ZN(G1342gat));
  AOI21_X1  g619(.A(G134gat), .B1(new_n799_), .B2(new_n580_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n552_), .A2(G134gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n808_), .B2(new_n822_), .ZN(G1343gat));
  AOI21_X1  g622(.A(new_n388_), .B1(new_n785_), .B2(new_n794_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n824_), .A2(new_n293_), .A3(new_n391_), .A4(new_n396_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n518_), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g626(.A1(new_n825_), .A2(new_n469_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT121), .B(G148gat), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1345gat));
  NOR2_X1   g629(.A1(new_n825_), .A2(new_n568_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT61), .B(G155gat), .Z(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1346gat));
  OR3_X1    g632(.A1(new_n825_), .A2(new_n537_), .A3(new_n621_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n537_), .B1(new_n825_), .B2(new_n549_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT122), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n834_), .A2(KEYINPUT122), .A3(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1347gat));
  NOR2_X1   g639(.A1(new_n396_), .A2(new_n293_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n388_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n612_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n805_), .A2(new_n667_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT123), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n805_), .A2(new_n846_), .A3(new_n667_), .A4(new_n843_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(G169gat), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT62), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n845_), .A2(new_n850_), .A3(G169gat), .A4(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n805_), .A2(new_n843_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT22), .B(G169gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n667_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT124), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n852_), .A2(new_n858_), .A3(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1348gat));
  AOI21_X1  g659(.A(G176gat), .B1(new_n853_), .B2(new_n470_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n391_), .B1(new_n785_), .B2(new_n794_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT125), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(G176gat), .A3(new_n470_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n842_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n861_), .B1(new_n865_), .B2(new_n866_), .ZN(G1349gat));
  NAND3_X1  g666(.A1(new_n863_), .A2(new_n633_), .A3(new_n866_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n567_), .A2(new_n294_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n868_), .A2(new_n561_), .B1(new_n853_), .B2(new_n869_), .ZN(G1350gat));
  NAND2_X1  g669(.A1(new_n853_), .A2(new_n552_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G190gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n853_), .A2(new_n580_), .A3(new_n295_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1351gat));
  NAND3_X1  g673(.A1(new_n824_), .A2(new_n391_), .A3(new_n841_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT126), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT126), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n824_), .A2(new_n877_), .A3(new_n391_), .A4(new_n841_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n518_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n513_), .ZN(G1352gat));
  AOI21_X1  g679(.A(new_n469_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT127), .B(G204gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1353gat));
  XNOR2_X1  g682(.A(KEYINPUT63), .B(G211gat), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n567_), .B(new_n884_), .C1(new_n876_), .C2(new_n878_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n876_), .A2(new_n878_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n588_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n885_), .B1(new_n887_), .B2(new_n888_), .ZN(G1354gat));
  AOI21_X1  g688(.A(G218gat), .B1(new_n886_), .B2(new_n580_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n621_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(G218gat), .B2(new_n891_), .ZN(G1355gat));
endmodule


