//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_;
  AND3_X1   g000(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n202_));
  AOI21_X1  g001(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT1), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT80), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n204_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n212_), .A2(new_n213_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n207_), .A2(new_n209_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n214_), .B(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n213_), .B(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n211_), .B(new_n217_), .C1(new_n219_), .C2(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n216_), .A2(KEYINPUT81), .A3(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT81), .B1(new_n216_), .B2(new_n222_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT4), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G127gat), .B(G134gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G113gat), .B(G120gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT79), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n216_), .A2(new_n229_), .A3(new_n222_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT4), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT91), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT92), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n231_), .A2(new_n234_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G1gat), .B(G29gat), .ZN(new_n242_));
  INV_X1    g041(.A(G85gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT0), .B(G57gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  NOR2_X1   g045(.A1(new_n241_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n246_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G197gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(G204gat), .ZN(new_n253_));
  INV_X1    g052(.A(G204gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n254_), .A2(G197gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT21), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(G197gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(G204gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT21), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n256_), .A2(new_n257_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT85), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT86), .B1(new_n253_), .B2(new_n255_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n257_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT86), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n258_), .A2(new_n259_), .A3(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n264_), .A2(new_n265_), .A3(KEYINPUT21), .A4(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT85), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n256_), .A2(new_n269_), .A3(new_n257_), .A4(new_n261_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n263_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT23), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(G183gat), .A3(G190gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT23), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT76), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n274_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT89), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n285_), .A2(KEYINPUT88), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT88), .B1(new_n285_), .B2(new_n286_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n284_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n275_), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT76), .B1(new_n275_), .B2(KEYINPUT23), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n273_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT89), .ZN(new_n293_));
  INV_X1    g092(.A(new_n281_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n282_), .A2(new_n283_), .A3(new_n289_), .A4(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G169gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(new_n284_), .A3(KEYINPUT75), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(G169gat), .B2(G176gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT24), .A3(new_n283_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n276_), .A2(new_n273_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT25), .B(G183gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT26), .B(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(new_n297_), .A3(new_n284_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n271_), .A2(new_n296_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT90), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT90), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n271_), .A2(new_n296_), .A3(new_n312_), .A4(new_n309_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT20), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n263_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n298_), .A2(new_n300_), .A3(new_n307_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n302_), .A2(new_n292_), .A3(new_n306_), .A4(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n303_), .A2(new_n294_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n285_), .A2(new_n286_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n284_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n320_), .A3(new_n283_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n314_), .B1(new_n315_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n311_), .A2(new_n313_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT19), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n296_), .A2(new_n309_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n315_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n315_), .A2(new_n322_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n330_), .A2(KEYINPUT20), .A3(new_n326_), .A4(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G8gat), .B(G36gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(G92gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT18), .B(G64gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n335_), .B(new_n336_), .Z(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n330_), .A2(KEYINPUT20), .A3(new_n327_), .A4(new_n331_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n310_), .A2(new_n323_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n326_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n337_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT94), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n337_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT94), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n338_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT27), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT27), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n328_), .A2(new_n343_), .A3(new_n332_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n338_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n251_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT29), .B1(new_n223_), .B2(new_n224_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT84), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n271_), .B1(G228gat), .B2(G233gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n358_), .B(KEYINPUT29), .C1(new_n223_), .C2(new_n224_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G78gat), .B(G106gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n216_), .B2(new_n222_), .ZN(new_n363_));
  OAI211_X1 g162(.A(G228gat), .B(G233gat), .C1(new_n271_), .C2(new_n363_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n360_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT87), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n360_), .A2(new_n364_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n361_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT87), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n360_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(G50gat), .B1(new_n225_), .B2(KEYINPUT29), .ZN(new_n374_));
  OR4_X1    g173(.A1(KEYINPUT29), .A2(new_n223_), .A3(new_n224_), .A4(G50gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT82), .B(G22gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT83), .B(KEYINPUT28), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n375_), .A3(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n367_), .A2(new_n373_), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n322_), .B(KEYINPUT30), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT78), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G15gat), .B(G43gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT77), .ZN(new_n388_));
  XOR2_X1   g187(.A(G71gat), .B(G99gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  XNOR2_X1  g191(.A(new_n322_), .B(KEYINPUT30), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT78), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n386_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n230_), .B(KEYINPUT31), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n390_), .B(new_n391_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT78), .A3(new_n385_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n396_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n397_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n380_), .A2(new_n382_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n403_), .B(KEYINPUT87), .C1(new_n365_), .C2(new_n366_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n384_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n402_), .B1(new_n384_), .B2(new_n404_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n354_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT32), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n333_), .B1(new_n408_), .B2(new_n343_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n342_), .A2(KEYINPUT32), .A3(new_n337_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n409_), .B(new_n410_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n241_), .B2(new_n246_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n239_), .A2(new_n240_), .A3(new_n248_), .A4(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n413_), .A2(new_n338_), .A3(new_n352_), .A4(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n231_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n232_), .A2(new_n233_), .A3(new_n238_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n246_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n411_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n384_), .A2(new_n404_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n402_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n407_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G230gat), .ZN(new_n425_));
  INV_X1    g224(.A(G233gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OAI22_X1  g229(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT65), .B1(KEYINPUT66), .B2(KEYINPUT7), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI221_X1 g232(.A(KEYINPUT65), .B1(KEYINPUT66), .B2(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT67), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n430_), .A2(new_n433_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G85gat), .B(G92gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n430_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT8), .B1(new_n440_), .B2(KEYINPUT67), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT68), .B1(new_n428_), .B2(new_n429_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G99gat), .A2(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT68), .ZN(new_n447_));
  NAND3_X1  g246(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n433_), .A2(new_n434_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n438_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT8), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n442_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT9), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n430_), .B1(new_n455_), .B2(new_n437_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT10), .B(G99gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT64), .ZN(new_n458_));
  INV_X1    g257(.A(G106gat), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n456_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(KEYINPUT9), .B2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G57gat), .B(G64gat), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n463_), .A2(KEYINPUT11), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(KEYINPUT11), .ZN(new_n465_));
  XOR2_X1   g264(.A(G71gat), .B(G78gat), .Z(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n465_), .A2(new_n466_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n454_), .A2(new_n462_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n439_), .A2(new_n441_), .B1(new_n452_), .B2(KEYINPUT8), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n461_), .A2(KEYINPUT9), .ZN(new_n473_));
  AOI211_X1 g272(.A(new_n473_), .B(new_n456_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n471_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(new_n475_), .A3(KEYINPUT12), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT12), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n477_), .B(new_n471_), .C1(new_n472_), .C2(new_n474_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n427_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT69), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n470_), .A2(new_n475_), .A3(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n482_), .B(new_n427_), .C1(new_n481_), .C2(new_n475_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G176gat), .B(G204gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G120gat), .B(G148gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n480_), .A2(new_n483_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT13), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n490_), .A2(KEYINPUT13), .A3(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G36gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G29gat), .ZN(new_n499_));
  INV_X1    g298(.A(G29gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G36gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT71), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n502_), .A2(KEYINPUT72), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT72), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(KEYINPUT71), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n499_), .B(new_n501_), .C1(new_n503_), .C2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n499_), .A2(new_n501_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n506_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516_));
  INV_X1    g315(.A(G1gat), .ZN(new_n517_));
  INV_X1    g316(.A(G8gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G1gat), .B(G8gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n515_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n522_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528_));
  INV_X1    g327(.A(new_n514_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n511_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n513_), .A2(KEYINPUT15), .A3(new_n514_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n527_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n515_), .A2(new_n522_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n533_), .A2(new_n525_), .A3(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G113gat), .B(G141gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G169gat), .B(G197gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  OR3_X1    g337(.A1(new_n526_), .A2(new_n535_), .A3(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n538_), .B1(new_n526_), .B2(new_n535_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n497_), .A2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n424_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G162gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT74), .B(G134gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n472_), .A2(new_n474_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n515_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n529_), .A2(new_n530_), .A3(new_n528_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT15), .B1(new_n513_), .B2(new_n514_), .ZN(new_n554_));
  OAI22_X1  g353(.A1(new_n472_), .A2(new_n474_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT34), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(KEYINPUT35), .A3(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(KEYINPUT35), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n556_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n566_), .A2(new_n560_), .B1(new_n555_), .B2(new_n552_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n545_), .B(new_n549_), .C1(new_n564_), .C2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n556_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n560_), .ZN(new_n570_));
  AOI211_X1 g369(.A(new_n565_), .B(new_n570_), .C1(new_n555_), .C2(new_n557_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n571_), .B2(new_n562_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n549_), .A2(new_n545_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n549_), .A2(new_n545_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n561_), .A2(new_n556_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n568_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT37), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n568_), .A2(new_n576_), .A3(KEYINPUT37), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n527_), .B(new_n469_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT17), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G127gat), .B(G155gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(G211gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(KEYINPUT16), .B(G183gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  OR3_X1    g389(.A1(new_n585_), .A2(new_n586_), .A3(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(KEYINPUT17), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n581_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n544_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT95), .Z(new_n597_));
  AND3_X1   g396(.A1(new_n597_), .A2(new_n517_), .A3(new_n251_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n598_), .A2(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n601_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n577_), .B(KEYINPUT97), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n594_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n544_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n250_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .A4(new_n610_), .ZN(G1324gat));
  AOI22_X1  g410(.A1(new_n333_), .A2(new_n337_), .B1(new_n347_), .B2(new_n346_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n351_), .B1(new_n612_), .B2(new_n345_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n353_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n518_), .B1(new_n608_), .B2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT39), .ZN(new_n617_));
  INV_X1    g416(.A(new_n615_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(G8gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n597_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g420(.A(G15gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n402_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n608_), .B2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n622_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n626_), .B1(new_n596_), .B2(new_n627_), .ZN(G1326gat));
  INV_X1    g427(.A(G22gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n422_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n608_), .B2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT42), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n629_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT100), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n632_), .B1(new_n596_), .B2(new_n634_), .ZN(G1327gat));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n568_), .A2(new_n576_), .A3(KEYINPUT37), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT37), .B1(new_n568_), .B2(new_n576_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT103), .B1(new_n424_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642_));
  AOI211_X1 g441(.A(new_n642_), .B(new_n639_), .C1(new_n407_), .C2(new_n423_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n579_), .A2(KEYINPUT102), .A3(new_n580_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n250_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n422_), .A2(new_n623_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n384_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n421_), .A2(new_n402_), .A3(new_n422_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n648_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT43), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n644_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n543_), .A2(new_n594_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT101), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n656_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(KEYINPUT44), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(KEYINPUT44), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n663_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n665_), .A2(new_n500_), .A3(new_n250_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n577_), .ZN(new_n667_));
  AND4_X1   g466(.A1(new_n667_), .A2(new_n424_), .A3(new_n594_), .A4(new_n543_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT105), .Z(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n251_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n666_), .A2(new_n670_), .ZN(G1328gat));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n498_), .A3(new_n615_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT45), .ZN(new_n673_));
  OAI21_X1  g472(.A(G36gat), .B1(new_n665_), .B2(new_n618_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(KEYINPUT46), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n675_), .B(new_n677_), .ZN(G1329gat));
  NAND3_X1  g477(.A1(new_n662_), .A2(new_n623_), .A3(new_n664_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n402_), .A2(G43gat), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n679_), .A2(G43gat), .B1(new_n669_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g481(.A(G50gat), .B1(new_n665_), .B2(new_n422_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n422_), .A2(G50gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT107), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n669_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(G1331gat));
  INV_X1    g486(.A(new_n497_), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n541_), .B(new_n688_), .C1(new_n407_), .C2(new_n423_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(new_n595_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n251_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n689_), .A2(new_n607_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n251_), .A2(G57gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(G1332gat));
  INV_X1    g493(.A(G64gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n692_), .B2(new_n615_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n615_), .A2(new_n695_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT109), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n690_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(G1333gat));
  INV_X1    g501(.A(G71gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n692_), .B2(new_n623_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT110), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT49), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n690_), .A2(new_n703_), .A3(new_n623_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1334gat));
  INV_X1    g507(.A(G78gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n692_), .B2(new_n630_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT50), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n690_), .A2(new_n709_), .A3(new_n630_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1335gat));
  INV_X1    g512(.A(new_n594_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n688_), .A2(new_n714_), .A3(new_n541_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n424_), .A3(new_n667_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n243_), .B1(new_n716_), .B2(new_n250_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT111), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n715_), .B(KEYINPUT113), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT112), .B1(new_n644_), .B2(new_n655_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n640_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n642_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n424_), .A2(KEYINPUT103), .A3(new_n640_), .ZN(new_n723_));
  AND4_X1   g522(.A1(KEYINPUT112), .A2(new_n655_), .A3(new_n722_), .A4(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n719_), .B1(new_n720_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT114), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT114), .B(new_n719_), .C1(new_n720_), .C2(new_n724_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n250_), .A2(new_n243_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n718_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT115), .Z(G1336gat));
  INV_X1    g531(.A(new_n716_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G92gat), .B1(new_n733_), .B2(new_n615_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n615_), .A2(G92gat), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT116), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n729_), .B2(new_n736_), .ZN(G1337gat));
  NAND3_X1  g536(.A1(new_n733_), .A2(new_n458_), .A3(new_n623_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n727_), .A2(new_n623_), .A3(new_n728_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n739_), .A2(KEYINPUT117), .A3(G99gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT117), .B1(new_n739_), .B2(G99gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n738_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT51), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(new_n738_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1338gat));
  NOR2_X1   g545(.A1(new_n656_), .A2(new_n422_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n459_), .B1(new_n747_), .B2(new_n719_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT52), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n733_), .A2(new_n459_), .A3(new_n630_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT53), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n749_), .A2(new_n753_), .A3(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1339gat));
  NOR2_X1   g554(.A1(new_n615_), .A2(new_n250_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n476_), .A2(new_n427_), .A3(new_n478_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT120), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(KEYINPUT55), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(KEYINPUT55), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n479_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n757_), .A2(KEYINPUT55), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT120), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n757_), .A2(new_n758_), .A3(KEYINPUT55), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n480_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n489_), .B1(new_n761_), .B2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n479_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n763_), .A2(new_n480_), .A3(new_n764_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n491_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT121), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n492_), .A2(new_n541_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT119), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n767_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n523_), .A2(new_n524_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n533_), .A2(new_n534_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT122), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n538_), .B(new_n777_), .C1(new_n779_), .C2(new_n524_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n493_), .A2(new_n539_), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n667_), .B1(new_n776_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT123), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n782_), .A2(new_n783_), .A3(KEYINPUT57), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n782_), .B2(KEYINPUT57), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n780_), .A2(new_n539_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n771_), .B2(new_n768_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n766_), .A2(KEYINPUT56), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n492_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n788_), .A2(new_n789_), .A3(KEYINPUT58), .A4(new_n492_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n776_), .A2(new_n781_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n577_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n794_), .A2(new_n581_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n714_), .B1(new_n786_), .B2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n595_), .A2(new_n542_), .A3(new_n688_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n801_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(KEYINPUT54), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n800_), .A2(new_n801_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n406_), .B(new_n756_), .C1(new_n799_), .C2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G113gat), .B1(new_n809_), .B2(new_n541_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT123), .B1(new_n796_), .B2(new_n797_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n796_), .A2(new_n797_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n792_), .A2(new_n793_), .A3(new_n581_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n782_), .A2(new_n783_), .A3(KEYINPUT57), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n594_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n807_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n650_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(KEYINPUT59), .A3(new_n756_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n542_), .B1(new_n812_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n810_), .B1(new_n822_), .B2(G113gat), .ZN(G1340gat));
  NOR2_X1   g622(.A1(new_n688_), .A2(G120gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n809_), .B1(KEYINPUT60), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n812_), .A2(new_n821_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n497_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G120gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(KEYINPUT60), .B2(new_n825_), .ZN(G1341gat));
  AOI21_X1  g628(.A(G127gat), .B1(new_n809_), .B2(new_n714_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n594_), .B1(new_n812_), .B2(new_n821_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g631(.A(G134gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n809_), .A2(new_n833_), .A3(new_n606_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n637_), .A2(new_n638_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n812_), .B2(new_n821_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n836_), .B2(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT124), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(new_n834_), .C1(new_n836_), .C2(new_n833_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1343gat));
  AOI21_X1  g640(.A(new_n651_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(new_n756_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n541_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n497_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT125), .B(G148gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1345gat));
  NAND3_X1  g647(.A1(new_n842_), .A2(new_n714_), .A3(new_n756_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G155gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1346gat));
  AOI21_X1  g651(.A(G162gat), .B1(new_n843_), .B2(new_n606_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n648_), .A2(G162gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n843_), .B2(new_n854_), .ZN(G1347gat));
  NOR2_X1   g654(.A1(new_n618_), .A2(new_n251_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n820_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n542_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n287_), .A2(new_n288_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n297_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT62), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n861_), .A2(KEYINPUT62), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1348gat));
  NOR2_X1   g663(.A1(new_n857_), .A2(new_n688_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n284_), .ZN(G1349gat));
  NOR2_X1   g665(.A1(new_n857_), .A2(new_n594_), .ZN(new_n867_));
  MUX2_X1   g666(.A(G183gat), .B(new_n304_), .S(new_n867_), .Z(G1350gat));
  OAI21_X1  g667(.A(G190gat), .B1(new_n857_), .B2(new_n835_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n606_), .A2(new_n305_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n857_), .B2(new_n870_), .ZN(G1351gat));
  NAND2_X1  g670(.A1(new_n842_), .A2(new_n856_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n542_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n252_), .ZN(G1352gat));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n688_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n254_), .ZN(G1353gat));
  INV_X1    g675(.A(new_n872_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT127), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n879_));
  INV_X1    g678(.A(G211gat), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n877_), .A2(new_n878_), .A3(new_n714_), .A4(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n842_), .A2(new_n714_), .A3(new_n856_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT127), .B1(new_n885_), .B2(new_n881_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n883_), .A2(new_n884_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n884_), .B1(new_n883_), .B2(new_n886_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1354gat));
  AND3_X1   g688(.A1(new_n877_), .A2(G218gat), .A3(new_n581_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G218gat), .B1(new_n877_), .B2(new_n606_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1355gat));
endmodule


