//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_;
  INV_X1    g000(.A(KEYINPUT105), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G204gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT89), .B1(new_n206_), .B2(G197gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT89), .ZN(new_n208_));
  INV_X1    g007(.A(G197gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(G204gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n206_), .A2(G197gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT90), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n205_), .A2(new_n212_), .A3(KEYINPUT90), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n212_), .A2(KEYINPUT21), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n206_), .A2(G197gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n209_), .A2(G204gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(KEYINPUT88), .B(KEYINPUT21), .C1(new_n219_), .C2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT21), .B1(new_n219_), .B2(new_n220_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT88), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n218_), .A2(new_n203_), .A3(new_n221_), .A4(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n217_), .A2(new_n225_), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n226_), .A2(KEYINPUT87), .B1(G228gat), .B2(G233gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(G141gat), .B2(G148gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n234_), .B1(new_n235_), .B2(KEYINPUT1), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT85), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n234_), .A2(KEYINPUT1), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n233_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n235_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n234_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT86), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(KEYINPUT86), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249_));
  INV_X1    g048(.A(G141gat), .ZN(new_n250_));
  INV_X1    g049(.A(G148gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .A4(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n230_), .A2(KEYINPUT2), .A3(new_n231_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n243_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n241_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n226_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n227_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n259_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G22gat), .B(G50gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n264_), .B(KEYINPUT28), .Z(new_n265_));
  XNOR2_X1  g064(.A(new_n263_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G78gat), .B(G106gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT91), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(KEYINPUT92), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n262_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(new_n268_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n273_), .B(new_n261_), .C1(new_n266_), .C2(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT20), .ZN(new_n277_));
  OR2_X1    g076(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n278_), .A2(KEYINPUT26), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G183gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT25), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT25), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(G190gat), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n282_), .B(new_n284_), .C1(KEYINPUT26), .C2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT81), .B1(new_n280_), .B2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n278_), .A2(KEYINPUT26), .A3(new_n279_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT25), .B(G183gat), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n285_), .A2(KEYINPUT26), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .A4(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G169gat), .ZN(new_n294_));
  INV_X1    g093(.A(G176gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  OR3_X1    g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n297_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n299_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n293_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n278_), .A2(new_n279_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n304_), .B1(G183gat), .B2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(KEYINPUT82), .B(G176gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G169gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n296_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n277_), .B1(new_n314_), .B2(new_n226_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT19), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT93), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n283_), .A2(G183gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n281_), .A2(KEYINPUT25), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n320_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT26), .B(G190gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n282_), .A2(new_n284_), .A3(KEYINPUT93), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT94), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n299_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n326_), .B2(new_n299_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n305_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT95), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n305_), .A2(new_n302_), .A3(KEYINPUT95), .A4(new_n303_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n328_), .A2(new_n329_), .A3(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n304_), .B1(G183gat), .B2(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n312_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n335_), .A2(new_n226_), .A3(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n319_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n224_), .A2(new_n203_), .A3(new_n221_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n342_), .A2(new_n218_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n293_), .A2(new_n306_), .B1(new_n312_), .B2(new_n309_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n277_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n326_), .A2(new_n299_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n334_), .B1(new_n346_), .B2(KEYINPUT94), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n326_), .A2(new_n327_), .A3(new_n299_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n338_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n345_), .B1(new_n343_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT96), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n317_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n350_), .B2(new_n317_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n341_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G64gat), .B(G92gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n360_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n362_), .B(new_n341_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT104), .B(KEYINPUT27), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n350_), .A2(new_n317_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT100), .B1(new_n335_), .B2(new_n338_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n347_), .A2(new_n348_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT100), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(new_n337_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n343_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n318_), .B1(new_n372_), .B2(new_n315_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n367_), .B1(new_n373_), .B2(KEYINPUT101), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT101), .ZN(new_n375_));
  AOI211_X1 g174(.A(new_n375_), .B(new_n318_), .C1(new_n372_), .C2(new_n315_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n360_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n343_), .B1(new_n369_), .B2(new_n337_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT20), .B1(new_n314_), .B2(new_n226_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n317_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT96), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n340_), .B1(new_n382_), .B2(new_n352_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n378_), .B1(new_n383_), .B2(new_n362_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n377_), .A2(KEYINPUT103), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT103), .B1(new_n377_), .B2(new_n384_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n276_), .B(new_n366_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(G127gat), .B(G134gat), .Z(new_n388_));
  XOR2_X1   g187(.A(G113gat), .B(G120gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G15gat), .B(G43gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT31), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G71gat), .B(G99gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n344_), .A2(KEYINPUT30), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n344_), .A2(KEYINPUT30), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n396_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n396_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n397_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n393_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n400_), .A2(new_n403_), .A3(new_n393_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n391_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n406_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n408_), .A2(new_n404_), .A3(KEYINPUT83), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n390_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(new_n391_), .A3(new_n406_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT83), .B1(new_n408_), .B2(new_n404_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n390_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT102), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT0), .ZN(new_n418_));
  INV_X1    g217(.A(G57gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G85gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n413_), .B1(new_n241_), .B2(new_n257_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n234_), .B(new_n242_), .C1(new_n253_), .C2(new_n255_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n238_), .A2(new_n240_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n424_), .B(new_n390_), .C1(new_n425_), .C2(new_n233_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n426_), .A3(KEYINPUT4), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT98), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT98), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n423_), .A2(new_n426_), .A3(new_n429_), .A4(KEYINPUT4), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n423_), .A2(KEYINPUT4), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n423_), .A2(new_n426_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n434_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n422_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  AOI211_X1 g239(.A(new_n421_), .B(new_n440_), .C1(new_n433_), .C2(new_n435_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n416_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n431_), .B1(new_n427_), .B2(KEYINPUT98), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n434_), .B1(new_n443_), .B2(new_n430_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n421_), .B1(new_n444_), .B2(new_n440_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n436_), .A2(new_n422_), .A3(new_n438_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(KEYINPUT102), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n415_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n202_), .B1(new_n387_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n365_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT103), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n350_), .A2(new_n317_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n371_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n343_), .B1(new_n349_), .B2(new_n370_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n315_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n317_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n455_), .B1(new_n459_), .B2(new_n375_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n376_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n362_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n363_), .A2(KEYINPUT27), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n454_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n377_), .A2(new_n384_), .A3(KEYINPUT103), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n453_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n448_), .B1(new_n414_), .B2(new_n410_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n466_), .A2(KEYINPUT105), .A3(new_n467_), .A4(new_n276_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n428_), .A2(new_n432_), .A3(new_n434_), .A4(new_n430_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n437_), .A2(new_n434_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n421_), .A2(new_n470_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n469_), .A2(new_n471_), .A3(KEYINPUT99), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT99), .B1(new_n469_), .B2(new_n471_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n361_), .A2(new_n363_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n439_), .A2(KEYINPUT33), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT33), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n445_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n362_), .A2(KEYINPUT32), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n480_), .ZN(new_n482_));
  OAI22_X1  g281(.A1(new_n355_), .A2(new_n482_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n483_));
  OAI22_X1  g282(.A1(new_n475_), .A2(new_n479_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n276_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n442_), .A2(new_n275_), .A3(new_n447_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n486_), .B(new_n366_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n415_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n451_), .A2(new_n468_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G127gat), .B(G155gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT16), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G183gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(G211gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT17), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n495_), .B(KEYINPUT78), .Z(new_n496_));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497_));
  INV_X1    g296(.A(G1gat), .ZN(new_n498_));
  INV_X1    g297(.A(G8gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G1gat), .B(G8gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  AND2_X1   g302(.A1(G231gat), .A2(G233gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G71gat), .B(G78gat), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G64gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(G57gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n419_), .A2(G64gat), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT67), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT67), .B1(new_n510_), .B2(new_n511_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT11), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT67), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n419_), .A2(G64gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n509_), .A2(G57gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT11), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT67), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n508_), .B1(new_n514_), .B2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n519_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(new_n507_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n522_), .A2(new_n524_), .A3(KEYINPUT69), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT69), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT11), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n507_), .B1(new_n527_), .B2(new_n523_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n514_), .A2(new_n508_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n526_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n506_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n505_), .B1(new_n530_), .B2(new_n525_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n496_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n528_), .A2(new_n529_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n505_), .B(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n494_), .A2(KEYINPUT17), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n495_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G29gat), .B(G36gat), .Z(new_n540_));
  XOR2_X1   g339(.A(G43gat), .B(G50gat), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G29gat), .B(G36gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT15), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT9), .ZN(new_n548_));
  INV_X1    g347(.A(G85gat), .ZN(new_n549_));
  INV_X1    g348(.A(G92gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G85gat), .A2(G92gat), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n548_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT66), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n557_));
  INV_X1    g356(.A(new_n552_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n557_), .B(new_n554_), .C1(new_n560_), .C2(new_n548_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n563_));
  INV_X1    g362(.A(G106gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT65), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT6), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n563_), .A2(KEYINPUT65), .A3(new_n564_), .A4(new_n565_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n568_), .A2(new_n571_), .A3(new_n572_), .A4(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n575_));
  INV_X1    g374(.A(G99gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n564_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n577_), .A2(new_n571_), .A3(new_n572_), .A4(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT8), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n579_), .A2(new_n580_), .A3(new_n560_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n579_), .B2(new_n560_), .ZN(new_n582_));
  OAI22_X1  g381(.A1(new_n562_), .A2(new_n574_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n547_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT34), .Z(new_n586_));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT74), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n542_), .A2(new_n545_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n590_), .B1(new_n583_), .B2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n584_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n586_), .A2(new_n587_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(KEYINPUT75), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n594_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT75), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n597_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n599_), .B(new_n600_), .C1(new_n584_), .C2(new_n592_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(KEYINPUT36), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n605_), .B(KEYINPUT36), .Z(new_n608_));
  NAND3_X1  g407(.A1(new_n595_), .A2(new_n601_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT37), .B1(new_n607_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT76), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT76), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n613_), .B(KEYINPUT37), .C1(new_n607_), .C2(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n602_), .A2(new_n606_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n616_), .A3(new_n609_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT77), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT77), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n615_), .A2(new_n619_), .A3(new_n616_), .A4(new_n609_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n612_), .A2(new_n614_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n490_), .A2(new_n539_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT64), .Z(new_n624_));
  NOR2_X1   g423(.A1(new_n535_), .A2(new_n583_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n582_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n579_), .A2(new_n580_), .A3(new_n560_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n571_), .A2(new_n572_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n567_), .B2(new_n566_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n630_), .A2(new_n556_), .A3(new_n561_), .A4(new_n573_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n628_), .A2(new_n631_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n624_), .B1(new_n625_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT68), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT12), .B1(new_n535_), .B2(new_n583_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n535_), .A2(new_n583_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n624_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT12), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n525_), .B2(new_n530_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n637_), .A2(new_n638_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT68), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n643_), .B(new_n624_), .C1(new_n625_), .C2(new_n632_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n634_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n645_), .A2(KEYINPUT70), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT70), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n634_), .A2(new_n642_), .A3(new_n653_), .A4(new_n644_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n655_), .B1(KEYINPUT72), .B2(KEYINPUT13), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n652_), .A2(new_n654_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT73), .Z(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n503_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n547_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n591_), .A2(KEYINPUT79), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT79), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n546_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n503_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n663_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(G229gat), .A2(G233gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n667_), .B(new_n503_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(G113gat), .B(G141gat), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(G169gat), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(new_n209_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n674_), .B(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n661_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n622_), .A2(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n681_), .A2(G1gat), .A3(new_n449_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n683_));
  OR2_X1    g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n490_), .A2(new_n539_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n659_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n679_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n607_), .A2(new_n610_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n688_), .A2(KEYINPUT107), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(KEYINPUT107), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n685_), .A2(new_n687_), .A3(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G1gat), .B1(new_n693_), .B2(new_n449_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n682_), .A2(new_n683_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n684_), .A2(new_n694_), .A3(new_n695_), .ZN(G1324gat));
  INV_X1    g495(.A(new_n466_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n685_), .A2(new_n697_), .A3(new_n687_), .A4(new_n692_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT39), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(G8gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G8gat), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n499_), .ZN(new_n702_));
  OAI22_X1  g501(.A1(new_n700_), .A2(new_n701_), .B1(new_n681_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g503(.A1(new_n681_), .A2(G15gat), .A3(new_n489_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT108), .ZN(new_n706_));
  OAI21_X1  g505(.A(G15gat), .B1(new_n693_), .B2(new_n489_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT41), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n707_), .A2(KEYINPUT41), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(KEYINPUT108), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n706_), .A2(new_n708_), .A3(new_n709_), .A4(new_n710_), .ZN(G1326gat));
  OR3_X1    g510(.A1(new_n681_), .A2(G22gat), .A3(new_n276_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n693_), .A2(new_n276_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G22gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G22gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1327gat));
  INV_X1    g516(.A(new_n539_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n688_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n490_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(new_n687_), .ZN(new_n721_));
  INV_X1    g520(.A(G29gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n448_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n451_), .A2(new_n468_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n415_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n724_), .B(new_n621_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n621_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n490_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n687_), .A2(new_n539_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n730_), .A2(KEYINPUT44), .A3(new_n732_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n448_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT109), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G29gat), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n737_), .A2(KEYINPUT109), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n723_), .B1(new_n739_), .B2(new_n740_), .ZN(G1328gat));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  INV_X1    g541(.A(G36gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT44), .B1(new_n730_), .B2(new_n732_), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n734_), .B(new_n731_), .C1(new_n727_), .C2(new_n729_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n743_), .B1(new_n746_), .B2(new_n697_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n720_), .A2(new_n743_), .A3(new_n697_), .A4(new_n687_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT111), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n748_), .B(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n742_), .B1(new_n747_), .B2(new_n752_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n744_), .A2(new_n745_), .A3(new_n466_), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT46), .B(new_n751_), .C1(new_n754_), .C2(new_n743_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1329gat));
  AOI21_X1  g555(.A(G43gat), .B1(new_n721_), .B2(new_n415_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n415_), .A2(G43gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n746_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(G1330gat));
  INV_X1    g560(.A(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n746_), .B2(new_n275_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n721_), .A2(new_n762_), .A3(new_n275_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT112), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n744_), .A2(new_n745_), .A3(new_n276_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n767_), .B(new_n764_), .C1(new_n768_), .C2(new_n762_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(G1331gat));
  NOR2_X1   g569(.A1(new_n660_), .A2(new_n678_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n685_), .A2(new_n692_), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n419_), .B1(new_n773_), .B2(new_n448_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n659_), .A2(new_n678_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n622_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n449_), .A2(G57gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n774_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT113), .ZN(G1332gat));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n509_), .A3(new_n697_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G64gat), .B1(new_n772_), .B2(new_n466_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(KEYINPUT48), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(KEYINPUT48), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n782_), .B2(new_n783_), .ZN(G1333gat));
  INV_X1    g583(.A(G71gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n776_), .A2(new_n785_), .A3(new_n415_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G71gat), .B1(new_n772_), .B2(new_n489_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(KEYINPUT49), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(KEYINPUT49), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n786_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT114), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n786_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1334gat));
  INV_X1    g593(.A(G78gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n776_), .A2(new_n795_), .A3(new_n275_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G78gat), .B1(new_n772_), .B2(new_n276_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n797_), .A2(KEYINPUT115), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(KEYINPUT115), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(KEYINPUT50), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT50), .B1(new_n798_), .B2(new_n799_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n796_), .B1(new_n800_), .B2(new_n801_), .ZN(G1335gat));
  AND2_X1   g601(.A1(new_n720_), .A2(new_n771_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G85gat), .B1(new_n803_), .B2(new_n448_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT116), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n775_), .A2(new_n539_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n808_), .A2(new_n549_), .A3(new_n449_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n805_), .A2(new_n809_), .ZN(G1336gat));
  OAI21_X1  g609(.A(G92gat), .B1(new_n808_), .B2(new_n466_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n803_), .A2(new_n550_), .A3(new_n697_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(G1337gat));
  OAI21_X1  g612(.A(G99gat), .B1(new_n808_), .B2(new_n489_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n803_), .A2(new_n415_), .A3(new_n563_), .A4(new_n565_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818_));
  OAI21_X1  g617(.A(G106gat), .B1(new_n818_), .B2(KEYINPUT117), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n807_), .B2(new_n275_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(KEYINPUT117), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n803_), .A2(new_n564_), .A3(new_n275_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT53), .B1(new_n822_), .B2(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1339gat));
  NOR4_X1   g628(.A1(new_n621_), .A2(new_n686_), .A3(new_n539_), .A4(new_n678_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT54), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n645_), .A2(new_n651_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n669_), .A2(KEYINPUT119), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n663_), .A2(new_n668_), .A3(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n671_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n677_), .B1(new_n673_), .B2(new_n670_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n674_), .A2(new_n677_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n832_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n642_), .A2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n637_), .A2(new_n641_), .A3(KEYINPUT55), .A4(new_n638_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n637_), .A2(new_n641_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n624_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n841_), .A2(new_n842_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n841_), .A2(new_n844_), .A3(KEYINPUT118), .A4(new_n842_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n651_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT56), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n650_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(KEYINPUT56), .A3(new_n848_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n839_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n854_), .A2(KEYINPUT58), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n621_), .B1(new_n854_), .B2(KEYINPUT58), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n678_), .A2(new_n832_), .ZN(new_n857_));
  AND4_X1   g656(.A1(KEYINPUT56), .A2(new_n847_), .A3(new_n651_), .A4(new_n848_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT56), .B1(new_n852_), .B2(new_n848_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n655_), .A2(new_n861_), .A3(new_n838_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n655_), .B2(new_n838_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n688_), .B1(new_n860_), .B2(new_n864_), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n855_), .A2(new_n856_), .B1(new_n865_), .B2(KEYINPUT57), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n865_), .A2(KEYINPUT57), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n831_), .B1(new_n868_), .B2(new_n539_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n387_), .A2(new_n449_), .A3(new_n489_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(G113gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n678_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT59), .B1(new_n869_), .B2(new_n871_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n867_), .B1(new_n866_), .B2(KEYINPUT121), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  OAI221_X1 g676(.A(new_n877_), .B1(new_n865_), .B2(KEYINPUT57), .C1(new_n855_), .C2(new_n856_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n718_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n831_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n871_), .A2(KEYINPUT59), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n875_), .B(new_n678_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n874_), .B1(new_n883_), .B2(new_n873_), .ZN(G1340gat));
  XNOR2_X1  g683(.A(KEYINPUT122), .B(G120gat), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n885_), .A2(KEYINPUT60), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n659_), .B2(KEYINPUT60), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n872_), .A2(new_n886_), .A3(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT123), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n875_), .B(new_n661_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n885_), .B2(new_n891_), .ZN(G1341gat));
  INV_X1    g691(.A(G127gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n872_), .A2(new_n893_), .A3(new_n718_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n875_), .B(new_n718_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n896_), .B2(new_n893_), .ZN(G1342gat));
  OAI21_X1  g696(.A(new_n875_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n898_));
  OAI21_X1  g697(.A(G134gat), .B1(new_n898_), .B2(new_n728_), .ZN(new_n899_));
  INV_X1    g698(.A(G134gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n872_), .A2(new_n900_), .A3(new_n691_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(G1343gat));
  NOR2_X1   g701(.A1(new_n869_), .A2(new_n415_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n903_), .A2(new_n275_), .A3(new_n448_), .A4(new_n466_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n679_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT124), .B(G141gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1344gat));
  NOR2_X1   g706(.A1(new_n904_), .A2(new_n660_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n251_), .ZN(G1345gat));
  NOR2_X1   g708(.A1(new_n904_), .A2(new_n539_), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT61), .B(G155gat), .Z(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT125), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n910_), .B(new_n912_), .ZN(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n904_), .B2(new_n728_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n692_), .A2(G162gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n904_), .B2(new_n915_), .ZN(G1347gat));
  NOR2_X1   g715(.A1(new_n466_), .A2(new_n450_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n275_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n678_), .B(new_n919_), .C1(new_n879_), .C2(new_n831_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G169gat), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n920_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n924_));
  INV_X1    g723(.A(new_n311_), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n920_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n923_), .A2(new_n924_), .A3(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT126), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n923_), .A2(new_n926_), .A3(new_n929_), .A4(new_n924_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1348gat));
  NOR3_X1   g730(.A1(new_n880_), .A2(new_n275_), .A3(new_n918_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n686_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n869_), .A2(new_n275_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n918_), .A2(new_n660_), .A3(new_n295_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n933_), .A2(new_n310_), .B1(new_n934_), .B2(new_n935_), .ZN(G1349gat));
  NOR2_X1   g735(.A1(new_n918_), .A2(new_n539_), .ZN(new_n937_));
  AOI21_X1  g736(.A(G183gat), .B1(new_n934_), .B2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n539_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n932_), .B2(new_n939_), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n932_), .A2(new_n324_), .A3(new_n691_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n932_), .A2(new_n621_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n285_), .ZN(G1351gat));
  NOR3_X1   g742(.A1(new_n466_), .A2(new_n276_), .A3(new_n448_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n903_), .A2(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n679_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n209_), .ZN(G1352gat));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n660_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(new_n206_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT127), .B(G204gat), .Z(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n948_), .B2(new_n951_), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n903_), .A2(new_n718_), .A3(new_n944_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  AND2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n953_), .A2(new_n954_), .A3(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n956_), .B1(new_n953_), .B2(new_n954_), .ZN(G1354gat));
  OAI21_X1  g756(.A(G218gat), .B1(new_n945_), .B2(new_n728_), .ZN(new_n958_));
  OR2_X1    g757(.A1(new_n692_), .A2(G218gat), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n945_), .B2(new_n959_), .ZN(G1355gat));
endmodule


