//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_;
  AND2_X1   g000(.A1(G57gat), .A2(G64gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G57gat), .A2(G64gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT69), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G57gat), .ZN(new_n205_));
  INV_X1    g004(.A(G64gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT69), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G57gat), .A2(G64gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n204_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT11), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT70), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n204_), .A2(new_n210_), .A3(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G71gat), .B(G78gat), .Z(new_n216_));
  AND2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n211_), .A2(new_n218_), .A3(KEYINPUT11), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n216_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n218_), .B1(new_n211_), .B2(KEYINPUT11), .ZN(new_n222_));
  AOI211_X1 g021(.A(KEYINPUT70), .B(new_n214_), .C1(new_n204_), .C2(new_n210_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT6), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT6), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(G99gat), .A3(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT10), .B(G99gat), .Z(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT66), .B1(G85gat), .B2(G92gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n235_));
  MUX2_X1   g034(.A(KEYINPUT66), .B(new_n234_), .S(new_n235_), .Z(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT65), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n230_), .B(new_n233_), .C1(new_n236_), .C2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT8), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n230_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT7), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n243_), .B(KEYINPUT67), .C1(G99gat), .C2(G106gat), .ZN(new_n244_));
  INV_X1    g043(.A(G99gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n245_), .B(new_n232_), .C1(new_n246_), .C2(KEYINPUT7), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n243_), .A2(KEYINPUT67), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n244_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n227_), .A2(new_n229_), .A3(KEYINPUT68), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n242_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G85gat), .B(G92gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n240_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  AOI211_X1 g053(.A(KEYINPUT8), .B(new_n252_), .C1(new_n249_), .C2(new_n230_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n239_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OR3_X1    g055(.A1(new_n225_), .A2(new_n256_), .A3(KEYINPUT71), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n249_), .A2(new_n230_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n240_), .A3(new_n253_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n243_), .A2(KEYINPUT67), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n246_), .A2(KEYINPUT7), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n245_), .A4(new_n232_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n262_), .A2(new_n244_), .B1(new_n230_), .B2(new_n241_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n252_), .B1(new_n263_), .B2(new_n250_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n259_), .B1(new_n264_), .B2(new_n240_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n265_), .A2(new_n239_), .B1(new_n220_), .B2(new_n224_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT72), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n265_), .A2(new_n220_), .A3(new_n224_), .A4(new_n239_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT71), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n225_), .A2(new_n256_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n257_), .A2(new_n267_), .A3(new_n269_), .A4(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G230gat), .A2(G233gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT64), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT12), .B1(new_n225_), .B2(new_n256_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(new_n266_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT12), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n225_), .A2(new_n256_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n275_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G120gat), .B(G148gat), .ZN(new_n284_));
  INV_X1    g083(.A(G204gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G176gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n268_), .A2(new_n270_), .A3(KEYINPUT12), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n276_), .B1(new_n291_), .B2(new_n281_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(new_n276_), .B2(new_n273_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n293_), .A2(new_n288_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT13), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT13), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n300_));
  OR2_X1    g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT86), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT2), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n307_));
  OAI221_X1 g106(.A(new_n307_), .B1(KEYINPUT84), .B2(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(new_n310_), .B2(KEYINPUT85), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n306_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n312_));
  OAI22_X1  g111(.A1(new_n305_), .A2(KEYINPUT2), .B1(new_n307_), .B2(KEYINPUT3), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n303_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT83), .B1(new_n302_), .B2(KEYINPUT1), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(G155gat), .A4(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n302_), .A2(KEYINPUT1), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n315_), .A2(new_n318_), .A3(new_n301_), .A4(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n320_), .B(new_n304_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n314_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT29), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT21), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G197gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(G204gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n285_), .A2(G197gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT21), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G211gat), .B(G218gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n329_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G211gat), .B(G218gat), .Z(new_n336_));
  OAI211_X1 g135(.A(new_n336_), .B(KEYINPUT21), .C1(new_n331_), .C2(new_n332_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G228gat), .A2(G233gat), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n326_), .A2(new_n338_), .B1(KEYINPUT88), .B2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n325_), .A2(KEYINPUT29), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G78gat), .B(G106gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n341_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n343_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n300_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n347_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n300_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n345_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G22gat), .B(G50gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n339_), .A2(KEYINPUT88), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n348_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT24), .ZN(new_n359_));
  INV_X1    g158(.A(G169gat), .ZN(new_n360_));
  INV_X1    g159(.A(G176gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G183gat), .A2(G190gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n362_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n368_));
  AND2_X1   g167(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n369_));
  AND2_X1   g168(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n371_));
  OAI22_X1  g170(.A1(new_n368_), .A2(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n360_), .A2(new_n361_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G169gat), .A2(G176gat), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT24), .A4(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(KEYINPUT24), .ZN(new_n377_));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT79), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n367_), .A2(new_n372_), .A3(new_n376_), .A4(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G183gat), .ZN(new_n381_));
  INV_X1    g180(.A(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n365_), .A2(new_n383_), .A3(new_n366_), .ZN(new_n384_));
  AND2_X1   g183(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n361_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n387_), .A3(new_n375_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n380_), .A2(new_n335_), .A3(new_n337_), .A4(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n389_), .A2(KEYINPUT20), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n375_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(KEYINPUT89), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT89), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n365_), .A2(new_n383_), .A3(new_n393_), .A4(new_n366_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n391_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n368_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n397_));
  OR2_X1    g196(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n396_), .A2(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n362_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n377_), .A2(new_n378_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n338_), .B1(new_n395_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n390_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G226gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT19), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n409_));
  AND3_X1   g208(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n372_), .A2(new_n412_), .A3(new_n362_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n379_), .A2(new_n376_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n388_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n409_), .B1(new_n415_), .B2(new_n338_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n391_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n393_), .B1(new_n412_), .B2(new_n383_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n394_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n367_), .B(new_n372_), .C1(new_n378_), .C2(new_n377_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n420_), .A2(new_n335_), .A3(new_n337_), .A4(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n407_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n416_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n408_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G92gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT18), .B(G64gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n408_), .B2(new_n424_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  OR3_X1    g232(.A1(new_n425_), .A2(KEYINPUT101), .A3(new_n429_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT97), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n390_), .A2(new_n435_), .A3(new_n423_), .A4(new_n404_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n404_), .A2(KEYINPUT20), .A3(new_n423_), .A4(new_n389_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT97), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n416_), .A2(new_n422_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n407_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n429_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT101), .B1(new_n425_), .B2(new_n429_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n434_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  MUX2_X1   g243(.A(new_n433_), .B(new_n444_), .S(KEYINPUT27), .Z(new_n445_));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n415_), .B(new_n446_), .Z(new_n447_));
  XNOR2_X1  g246(.A(G127gat), .B(G134gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G113gat), .B(G120gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT31), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT81), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n447_), .B(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(KEYINPUT80), .B(G43gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT30), .B(G15gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n453_), .B(new_n458_), .Z(new_n459_));
  NAND3_X1  g258(.A1(new_n358_), .A2(new_n445_), .A3(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G1gat), .B(G29gat), .ZN(new_n461_));
  INV_X1    g260(.A(G85gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT0), .B(G57gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n314_), .A2(new_n324_), .A3(new_n450_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n450_), .B1(new_n314_), .B2(new_n324_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT90), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n471_));
  INV_X1    g270(.A(new_n450_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n325_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n467_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT92), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n325_), .A2(new_n472_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n314_), .A2(new_n324_), .A3(new_n450_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n471_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n325_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(KEYINPUT90), .A3(new_n450_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT92), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n467_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n475_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT91), .B(KEYINPUT4), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n476_), .A2(new_n485_), .ZN(new_n486_));
  AOI211_X1 g285(.A(new_n467_), .B(new_n486_), .C1(new_n481_), .C2(KEYINPUT4), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n466_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT4), .B1(new_n470_), .B2(new_n473_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n467_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n486_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n492_), .A2(new_n475_), .A3(new_n465_), .A4(new_n483_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n460_), .A2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT94), .B(KEYINPUT33), .Z(new_n496_));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n482_), .B1(new_n481_), .B2(new_n467_), .ZN(new_n499_));
  AOI211_X1 g298(.A(KEYINPUT92), .B(new_n490_), .C1(new_n478_), .C2(new_n480_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n501_), .A2(KEYINPUT93), .A3(new_n465_), .A4(new_n492_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n498_), .A2(KEYINPUT95), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT95), .B1(new_n498_), .B2(new_n502_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n501_), .A2(KEYINPUT33), .A3(new_n465_), .A4(new_n492_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n489_), .A2(new_n467_), .A3(new_n491_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n465_), .B1(new_n481_), .B2(new_n490_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT96), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n506_), .A2(KEYINPUT96), .A3(new_n507_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n505_), .B(new_n433_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n503_), .A2(new_n504_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n431_), .A2(KEYINPUT32), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n441_), .A2(KEYINPUT98), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT98), .B1(new_n441_), .B2(new_n513_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n408_), .A2(new_n424_), .A3(new_n512_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n494_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT99), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT99), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n465_), .B1(new_n501_), .B2(new_n492_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n493_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n517_), .B(new_n520_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n519_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n358_), .B1(new_n511_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT100), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n494_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n357_), .A2(new_n528_), .A3(new_n445_), .ZN(new_n529_));
  OAI211_X1 g328(.A(KEYINPUT100), .B(new_n358_), .C1(new_n511_), .C2(new_n524_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n459_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n495_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT76), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT75), .B(G1gat), .ZN(new_n535_));
  INV_X1    g334(.A(G8gat), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT14), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G1gat), .B(G8gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n541_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G29gat), .B(G36gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n547_), .A2(KEYINPUT15), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(KEYINPUT15), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n543_), .B(new_n544_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n544_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n547_), .B1(new_n551_), .B2(new_n542_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n534_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n551_), .A2(new_n542_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n547_), .B(KEYINPUT15), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT76), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n553_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n545_), .B(new_n546_), .Z(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n557_), .B1(new_n561_), .B2(new_n552_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G169gat), .B(G197gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT78), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT77), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n563_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT102), .B1(new_n533_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n530_), .A2(new_n529_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n523_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n520_), .B1(new_n494_), .B2(new_n517_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n493_), .A2(new_n497_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n496_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n502_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT95), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n498_), .A2(KEYINPUT95), .A3(new_n502_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n505_), .A2(new_n433_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n509_), .A2(new_n508_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n575_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT100), .B1(new_n586_), .B2(new_n358_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n532_), .B1(new_n572_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n495_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT102), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n569_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n299_), .B1(new_n571_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT34), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT35), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n256_), .B2(new_n555_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n265_), .A2(new_n239_), .A3(new_n547_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n597_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT74), .ZN(new_n603_));
  INV_X1    g402(.A(new_n598_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n601_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(KEYINPUT73), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n605_), .A2(KEYINPUT73), .B1(new_n256_), .B2(new_n555_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n604_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n603_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610_));
  XOR2_X1   g409(.A(G190gat), .B(G218gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n609_), .A2(new_n610_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n610_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n613_), .A2(new_n610_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n615_), .B(new_n616_), .C1(new_n603_), .C2(new_n608_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n614_), .A2(KEYINPUT37), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT37), .B1(new_n614_), .B2(new_n617_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n554_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(new_n225_), .ZN(new_n624_));
  XOR2_X1   g423(.A(G127gat), .B(G155gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(G211gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(KEYINPUT16), .B(G183gat), .Z(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT17), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n624_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n624_), .A2(KEYINPUT17), .A3(new_n628_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n621_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n593_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n494_), .A3(new_n535_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n638_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n299_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(KEYINPUT104), .A3(new_n569_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(new_n299_), .B2(new_n570_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n614_), .A2(new_n617_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n633_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n590_), .A2(new_n645_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G1gat), .B1(new_n650_), .B2(new_n528_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n639_), .A2(new_n640_), .A3(new_n651_), .ZN(G1324gat));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n653_));
  INV_X1    g452(.A(new_n445_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n649_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n656_), .B2(KEYINPUT39), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(KEYINPUT39), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n655_), .A2(KEYINPUT105), .A3(new_n659_), .A4(G8gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n635_), .A2(new_n536_), .A3(new_n654_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(new_n662_), .A3(KEYINPUT40), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1325gat));
  INV_X1    g466(.A(G15gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n649_), .B2(new_n459_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT41), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n635_), .A2(new_n668_), .A3(new_n459_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1326gat));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n649_), .B2(new_n357_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT42), .Z(new_n675_));
  NAND3_X1  g474(.A1(new_n635_), .A2(new_n673_), .A3(new_n357_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1327gat));
  NOR2_X1   g476(.A1(new_n646_), .A2(new_n632_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n592_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n591_), .B1(new_n590_), .B2(new_n569_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n641_), .B(new_n678_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n494_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n642_), .A2(new_n633_), .A3(new_n644_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT43), .B1(new_n533_), .B2(new_n620_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n590_), .A2(new_n688_), .A3(new_n621_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n686_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT108), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n686_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n688_), .B1(new_n590_), .B2(new_n621_), .ZN(new_n694_));
  AOI211_X1 g493(.A(KEYINPUT43), .B(new_n620_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697_));
  INV_X1    g496(.A(new_n691_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n696_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n690_), .A2(KEYINPUT44), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n692_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n494_), .A2(G29gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n683_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  NAND4_X1  g502(.A1(new_n692_), .A2(new_n699_), .A3(new_n654_), .A4(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G36gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n706_));
  NOR2_X1   g505(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n445_), .A2(G36gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT45), .B1(new_n681_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n593_), .A2(new_n711_), .A3(new_n678_), .A4(new_n708_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n705_), .A2(new_n706_), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n706_), .B1(new_n705_), .B2(new_n713_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1329gat));
  NAND3_X1  g515(.A1(new_n692_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n459_), .A2(G43gat), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n681_), .A2(new_n532_), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n717_), .A2(new_n718_), .B1(G43gat), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n717_), .B2(new_n358_), .ZN(new_n722_));
  INV_X1    g521(.A(G50gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n682_), .A2(new_n723_), .A3(new_n357_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n641_), .A2(new_n569_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n590_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n648_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n728_), .A2(new_n205_), .A3(new_n528_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n634_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n494_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n729_), .B1(new_n205_), .B2(new_n732_), .ZN(G1332gat));
  OAI21_X1  g532(.A(G64gat), .B1(new_n728_), .B2(new_n445_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n206_), .A3(new_n654_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(KEYINPUT110), .A3(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1333gat));
  OAI21_X1  g540(.A(G71gat), .B1(new_n728_), .B2(new_n532_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n532_), .A2(G71gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n730_), .B2(new_n745_), .ZN(G1334gat));
  OAI21_X1  g545(.A(G78gat), .B1(new_n728_), .B2(new_n358_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT50), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n358_), .A2(G78gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n730_), .B2(new_n749_), .ZN(G1335gat));
  NAND2_X1  g549(.A1(new_n727_), .A2(new_n678_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n494_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n726_), .A2(new_n633_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n528_), .A2(new_n462_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n755_), .B2(new_n756_), .ZN(G1336gat));
  AOI21_X1  g556(.A(G92gat), .B1(new_n752_), .B2(new_n654_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n654_), .A2(G92gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n755_), .B2(new_n759_), .ZN(G1337gat));
  AOI21_X1  g559(.A(new_n245_), .B1(new_n755_), .B2(new_n459_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n459_), .A2(new_n231_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n752_), .B2(new_n762_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g563(.A1(new_n752_), .A2(new_n232_), .A3(new_n357_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n755_), .A2(new_n357_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G106gat), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT52), .B(new_n232_), .C1(new_n755_), .C2(new_n357_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g570(.A1(new_n569_), .A2(G113gat), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT119), .Z(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n460_), .A2(new_n528_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n632_), .A2(new_n570_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT112), .Z(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n641_), .A3(new_n620_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n283_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n291_), .A2(new_n276_), .A3(new_n281_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n291_), .A2(KEYINPUT113), .A3(new_n276_), .A4(new_n281_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n292_), .A2(KEYINPUT55), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n784_), .A2(new_n787_), .A3(new_n788_), .A4(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n288_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n791_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n790_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n791_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n559_), .A2(new_n567_), .A3(new_n562_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n567_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n558_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n561_), .A2(new_n557_), .A3(new_n552_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n797_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n289_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n803_), .A2(KEYINPUT114), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(KEYINPUT114), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n795_), .A2(new_n796_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n621_), .B1(new_n806_), .B2(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n795_), .A2(new_n796_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n804_), .A2(new_n805_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(KEYINPUT58), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(KEYINPUT116), .A3(KEYINPUT58), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n807_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n569_), .A2(new_n289_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n793_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(new_n792_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n295_), .A2(new_n801_), .A3(new_n797_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n646_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n633_), .B1(new_n814_), .B2(new_n821_), .ZN(new_n822_));
  AOI211_X1 g621(.A(KEYINPUT59), .B(new_n776_), .C1(new_n782_), .C2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n808_), .A2(new_n809_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n620_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827_));
  AND4_X1   g626(.A1(KEYINPUT116), .A2(new_n808_), .A3(KEYINPUT58), .A4(new_n809_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT116), .B1(new_n806_), .B2(KEYINPUT58), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n826_), .B(new_n827_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n819_), .B(KEYINPUT57), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n812_), .A2(new_n813_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n827_), .B1(new_n833_), .B2(new_n826_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n633_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n776_), .B1(new_n835_), .B2(new_n782_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT118), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n826_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT117), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n781_), .B1(new_n842_), .B2(new_n633_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n839_), .B(KEYINPUT59), .C1(new_n843_), .C2(new_n776_), .ZN(new_n844_));
  AOI211_X1 g643(.A(new_n774_), .B(new_n823_), .C1(new_n838_), .C2(new_n844_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n843_), .A2(new_n570_), .A3(new_n776_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(G113gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT120), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n823_), .B1(new_n838_), .B2(new_n844_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n773_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851_));
  INV_X1    g650(.A(new_n847_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n848_), .A2(new_n853_), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n641_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n836_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n849_), .A2(new_n299_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n855_), .ZN(G1341gat));
  AOI21_X1  g658(.A(G127gat), .B1(new_n836_), .B2(new_n632_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n633_), .A2(KEYINPUT121), .ZN(new_n861_));
  MUX2_X1   g660(.A(KEYINPUT121), .B(new_n861_), .S(G127gat), .Z(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n849_), .B2(new_n862_), .ZN(G1342gat));
  AOI21_X1  g662(.A(G134gat), .B1(new_n836_), .B2(new_n647_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n621_), .A2(G134gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n849_), .B2(new_n865_), .ZN(G1343gat));
  NOR2_X1   g665(.A1(new_n358_), .A2(new_n654_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n494_), .A3(new_n532_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT122), .B1(new_n843_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n870_));
  INV_X1    g669(.A(new_n868_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n821_), .B1(new_n814_), .B2(new_n827_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n632_), .B1(new_n872_), .B2(new_n841_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n870_), .B(new_n871_), .C1(new_n873_), .C2(new_n781_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n869_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n569_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n299_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n875_), .B2(new_n632_), .ZN(new_n881_));
  AOI211_X1 g680(.A(KEYINPUT123), .B(new_n633_), .C1(new_n869_), .C2(new_n874_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n881_), .A2(new_n882_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n835_), .A2(new_n782_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n870_), .B1(new_n886_), .B2(new_n871_), .ZN(new_n887_));
  AOI211_X1 g686(.A(KEYINPUT122), .B(new_n868_), .C1(new_n835_), .C2(new_n782_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n632_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT123), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n875_), .A2(new_n880_), .A3(new_n632_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n883_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n885_), .A2(new_n892_), .ZN(G1346gat));
  AOI21_X1  g692(.A(G162gat), .B1(new_n875_), .B2(new_n647_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n621_), .A2(G162gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n875_), .B2(new_n895_), .ZN(G1347gat));
  NOR3_X1   g695(.A1(new_n445_), .A2(new_n494_), .A3(new_n532_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  AOI211_X1 g697(.A(new_n357_), .B(new_n898_), .C1(new_n782_), .C2(new_n822_), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n899_), .B(new_n569_), .C1(new_n386_), .C2(new_n385_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n360_), .B1(new_n899_), .B2(new_n569_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(KEYINPUT124), .A3(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n904_));
  AOI21_X1  g703(.A(KEYINPUT124), .B1(new_n901_), .B2(new_n902_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n900_), .B1(new_n904_), .B2(new_n905_), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n899_), .B2(new_n299_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n843_), .A2(new_n357_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n898_), .A2(new_n641_), .A3(new_n361_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n908_), .B2(new_n909_), .ZN(G1349gat));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n632_), .A3(new_n897_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n633_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n911_), .A2(new_n381_), .B1(new_n899_), .B2(new_n912_), .ZN(G1350gat));
  AOI21_X1  g712(.A(new_n382_), .B1(new_n899_), .B2(new_n621_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT125), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n899_), .B(new_n647_), .C1(new_n371_), .C2(new_n370_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1351gat));
  NOR4_X1   g716(.A1(new_n358_), .A2(new_n494_), .A3(new_n445_), .A4(new_n459_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n886_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n921_), .A2(new_n330_), .A3(new_n570_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n919_), .B(KEYINPUT126), .ZN(new_n923_));
  AOI21_X1  g722(.A(G197gat), .B1(new_n923_), .B2(new_n569_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1352gat));
  OAI211_X1 g724(.A(KEYINPUT127), .B(G204gat), .C1(new_n921_), .C2(new_n641_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n923_), .A2(new_n299_), .A3(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1353gat));
  XNOR2_X1  g728(.A(KEYINPUT63), .B(G211gat), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n921_), .A2(new_n633_), .A3(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n923_), .A2(new_n632_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n931_), .B1(new_n932_), .B2(new_n933_), .ZN(G1354gat));
  AND3_X1   g733(.A1(new_n923_), .A2(G218gat), .A3(new_n621_), .ZN(new_n935_));
  AOI21_X1  g734(.A(G218gat), .B1(new_n923_), .B2(new_n647_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1355gat));
endmodule


