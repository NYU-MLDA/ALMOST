//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G22gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G15gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G1gat), .B(G8gat), .Z(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n203_), .A2(new_n208_), .A3(new_n206_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n215_));
  XOR2_X1   g014(.A(G71gat), .B(G78gat), .Z(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n215_), .A2(new_n216_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n212_), .B(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G231gat), .A2(G233gat), .ZN(new_n221_));
  XOR2_X1   g020(.A(new_n220_), .B(new_n221_), .Z(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G183gat), .B(G211gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G127gat), .B(G155gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  OR3_X1    g028(.A1(new_n223_), .A2(new_n224_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(KEYINPUT17), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n223_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT37), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G190gat), .B(G218gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G134gat), .B(G162gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT36), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n239_), .A2(KEYINPUT69), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n239_), .A2(KEYINPUT69), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n244_));
  OR3_X1    g043(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT6), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT65), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT6), .ZN(new_n249_));
  AND2_X1   g048(.A1(G99gat), .A2(G106gat), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n247_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n244_), .B(new_n245_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT8), .ZN(new_n254_));
  XOR2_X1   g053(.A(G85gat), .B(G92gat), .Z(new_n255_));
  AND3_X1   g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT66), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT8), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(G85gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(G85gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(KEYINPUT9), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT10), .B(G99gat), .Z(new_n269_));
  INV_X1    g068(.A(G106gat), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n268_), .A2(G92gat), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n255_), .A2(KEYINPUT9), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n271_), .B(new_n272_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n264_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G29gat), .B(G36gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G43gat), .B(G50gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT15), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n273_), .B(new_n277_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G232gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT34), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n279_), .B(new_n280_), .C1(KEYINPUT35), .C2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(KEYINPUT35), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n283_), .A2(new_n285_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n241_), .B(new_n243_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n237_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(KEYINPUT36), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n292_), .A3(new_n286_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n234_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n239_), .B1(new_n290_), .B2(new_n286_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(new_n234_), .A3(new_n293_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n233_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT72), .ZN(new_n300_));
  INV_X1    g099(.A(new_n219_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n274_), .A2(KEYINPUT12), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G230gat), .A2(G233gat), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n273_), .B(new_n219_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT12), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n273_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n301_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n302_), .A2(new_n303_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n304_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n303_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G176gat), .B(G204gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G120gat), .B(G148gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n313_), .A2(new_n319_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n321_), .A2(new_n322_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n210_), .A2(new_n211_), .A3(new_n277_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n212_), .B2(new_n278_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G229gat), .A2(G233gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n330_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n212_), .A2(new_n278_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT73), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n277_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n339_));
  OAI211_X1 g138(.A(G229gat), .B(G233gat), .C1(new_n330_), .C2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n334_), .A2(new_n338_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G113gat), .B(G141gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G169gat), .B(G197gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(KEYINPUT74), .A3(new_n344_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n344_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n334_), .A2(new_n338_), .A3(new_n340_), .A4(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT75), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355_));
  INV_X1    g154(.A(G169gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT77), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(G169gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n359_), .A3(KEYINPUT22), .ZN(new_n360_));
  INV_X1    g159(.A(G176gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n363_));
  NOR2_X1   g162(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n364_));
  OAI21_X1  g163(.A(G169gat), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT79), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n367_), .B(G169gat), .C1(new_n363_), .C2(new_n364_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n362_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n355_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT23), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(G183gat), .B2(G190gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT77), .B(G169gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(G176gat), .B1(new_n376_), .B2(KEYINPUT22), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT78), .B(KEYINPUT22), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n367_), .B1(new_n378_), .B2(G169gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n368_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n377_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(KEYINPUT80), .A3(new_n370_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n372_), .A2(new_n375_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n356_), .A2(new_n361_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n385_), .A2(KEYINPUT24), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(KEYINPUT24), .A3(new_n370_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n374_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT76), .B1(new_n390_), .B2(G183gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT25), .B(G183gat), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n389_), .B(new_n391_), .C1(new_n392_), .C2(KEYINPUT76), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n383_), .A2(new_n384_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n384_), .B1(new_n383_), .B2(new_n394_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT81), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n383_), .A2(new_n394_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT30), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n383_), .A2(new_n384_), .A3(new_n394_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G15gat), .B(G43gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G99gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405_));
  INV_X1    g204(.A(G71gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n404_), .B(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n397_), .A2(new_n402_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n408_), .ZN(new_n410_));
  OAI211_X1 g209(.A(KEYINPUT81), .B(new_n410_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n409_), .A2(KEYINPUT83), .A3(new_n411_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416_));
  OR2_X1    g215(.A1(G127gat), .A2(G134gat), .ZN(new_n417_));
  INV_X1    g216(.A(G120gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G113gat), .ZN(new_n419_));
  INV_X1    g218(.A(G113gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G120gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G127gat), .A2(G134gat), .ZN(new_n422_));
  AND4_X1   g221(.A1(new_n417_), .A2(new_n419_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n419_), .A2(new_n421_), .B1(new_n417_), .B2(new_n422_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n416_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n417_), .A2(new_n422_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n419_), .A2(new_n421_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n417_), .A2(new_n419_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(KEYINPUT82), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n431_), .B(KEYINPUT31), .Z(new_n432_));
  NAND3_X1  g231(.A1(new_n414_), .A2(new_n415_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT1), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(G155gat), .B2(G162gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G155gat), .A2(G162gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT84), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(G155gat), .A3(G162gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n436_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G155gat), .A2(G162gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT1), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n437_), .A2(new_n438_), .A3(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(G141gat), .B(G148gat), .Z(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n423_), .A2(new_n424_), .ZN(new_n447_));
  OR3_X1    g246(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G141gat), .A2(G148gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT2), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n448_), .A2(new_n451_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n440_), .A3(new_n439_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n446_), .A2(new_n447_), .A3(new_n455_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n446_), .A2(new_n455_), .B1(new_n425_), .B2(new_n430_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT89), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n454_), .A2(new_n439_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n459_), .A2(new_n440_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n447_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n458_), .A2(KEYINPUT4), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT90), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G225gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n446_), .A2(new_n455_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n431_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n469_), .A2(KEYINPUT4), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n458_), .A2(new_n463_), .A3(new_n471_), .A4(KEYINPUT4), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n465_), .A2(new_n467_), .A3(new_n470_), .A4(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n458_), .A2(new_n466_), .A3(new_n463_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G85gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G29gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  AND3_X1   g278(.A1(new_n473_), .A2(new_n474_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n432_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n409_), .A2(KEYINPUT83), .A3(new_n411_), .A4(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n433_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT93), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT29), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n460_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT28), .B(G22gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(G50gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n488_), .B(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G78gat), .B(G106gat), .Z(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G197gat), .B(G204gat), .ZN(new_n494_));
  AND2_X1   g293(.A1(G211gat), .A2(G218gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(G211gat), .A2(G218gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT21), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n494_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(G211gat), .A2(G218gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G211gat), .A2(G218gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G197gat), .B(G204gat), .Z(new_n504_));
  NAND3_X1  g303(.A1(new_n501_), .A2(KEYINPUT86), .A3(new_n502_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT21), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n500_), .A2(KEYINPUT85), .A3(new_n503_), .A4(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G228gat), .A2(G233gat), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n487_), .B1(new_n446_), .B2(new_n455_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n500_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n509_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n508_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n511_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n513_), .B(new_n514_), .C1(new_n460_), .C2(new_n487_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n493_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n491_), .B1(new_n516_), .B2(KEYINPUT87), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT88), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n491_), .B(new_n519_), .C1(new_n516_), .C2(KEYINPUT87), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n516_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n512_), .A2(new_n515_), .A3(new_n493_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n518_), .A2(new_n522_), .A3(new_n523_), .A4(new_n520_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G8gat), .B(G36gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G92gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT18), .B(G64gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  NAND2_X1  g330(.A1(G226gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT19), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT20), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n398_), .B2(new_n514_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n392_), .A2(new_n389_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n388_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT22), .B(G169gat), .Z(new_n538_));
  OAI21_X1  g337(.A(new_n375_), .B1(G176gat), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n539_), .B2(new_n371_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(new_n514_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n533_), .B1(new_n535_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n383_), .A2(new_n511_), .A3(new_n394_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n514_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n544_), .A2(KEYINPUT20), .A3(new_n533_), .A4(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n531_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n531_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n533_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n535_), .B2(new_n542_), .ZN(new_n551_));
  AND4_X1   g350(.A1(KEYINPUT20), .A2(new_n544_), .A3(new_n550_), .A4(new_n545_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n549_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n548_), .A2(new_n553_), .A3(KEYINPUT27), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n535_), .A2(new_n542_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n550_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT27), .B1(new_n557_), .B2(new_n548_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n527_), .A2(new_n554_), .A3(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n485_), .A2(new_n486_), .A3(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n433_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT27), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n549_), .B1(new_n556_), .B2(new_n546_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n543_), .A2(new_n547_), .A3(new_n531_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n548_), .A2(new_n553_), .A3(KEYINPUT27), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n565_), .A2(new_n526_), .A3(new_n525_), .A4(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT93), .B1(new_n561_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n560_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n433_), .A2(new_n484_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n563_), .A2(new_n564_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n473_), .A2(KEYINPUT33), .A3(new_n474_), .A4(new_n479_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n462_), .B1(new_n461_), .B2(new_n469_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n456_), .A2(KEYINPUT89), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT92), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n458_), .A2(new_n577_), .A3(new_n463_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n467_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n479_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n465_), .A2(new_n466_), .A3(new_n470_), .A4(new_n472_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n573_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n571_), .B(new_n572_), .C1(new_n583_), .C2(new_n480_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n531_), .A2(KEYINPUT32), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n586_));
  OAI211_X1 g385(.A(KEYINPUT32), .B(new_n531_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n586_), .B(new_n587_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n527_), .B1(new_n584_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n482_), .A2(new_n527_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n565_), .A2(new_n566_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n570_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n593_));
  AOI211_X1 g392(.A(new_n329_), .B(new_n354_), .C1(new_n569_), .C2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n300_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT94), .ZN(new_n596_));
  INV_X1    g395(.A(new_n482_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n204_), .A3(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n290_), .A2(new_n292_), .A3(new_n286_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(new_n296_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(new_n233_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n594_), .A2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n604_), .A2(new_n597_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n600_), .B1(new_n204_), .B2(new_n605_), .ZN(G1324gat));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n591_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n607_), .A2(G8gat), .B1(KEYINPUT96), .B2(new_n608_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n609_), .A2(KEYINPUT96), .A3(new_n608_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n596_), .A2(new_n205_), .A3(new_n591_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(KEYINPUT96), .B2(new_n608_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT40), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(G1325gat));
  INV_X1    g414(.A(new_n570_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n604_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(G15gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT41), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n595_), .A2(G15gat), .A3(new_n570_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1326gat));
  NAND2_X1  g420(.A1(new_n604_), .A2(new_n527_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G22gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT42), .ZN(new_n624_));
  INV_X1    g423(.A(new_n527_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n625_), .A2(G22gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n595_), .B2(new_n626_), .ZN(G1327gat));
  NAND2_X1  g426(.A1(new_n569_), .A2(new_n593_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n233_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n329_), .A2(new_n629_), .A3(new_n354_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n628_), .A2(new_n602_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(G29gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(new_n597_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n295_), .A2(new_n298_), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT43), .B(new_n634_), .C1(new_n569_), .C2(new_n593_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n569_), .A2(new_n593_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n569_), .B2(new_n593_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n295_), .A2(new_n640_), .A3(new_n298_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n601_), .A2(new_n296_), .A3(KEYINPUT37), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT99), .B1(new_n642_), .B2(new_n294_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n638_), .A2(new_n639_), .A3(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT97), .B(KEYINPUT43), .Z(new_n646_));
  OAI21_X1  g445(.A(new_n636_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n630_), .B1(new_n648_), .B2(KEYINPUT44), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(KEYINPUT44), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n647_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n651_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n486_), .B1(new_n485_), .B2(new_n559_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n561_), .A2(new_n567_), .A3(KEYINPUT93), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n473_), .A2(new_n474_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n582_), .A2(new_n580_), .A3(new_n579_), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n657_), .A2(new_n479_), .B1(new_n658_), .B2(KEYINPUT33), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n572_), .A2(new_n548_), .A3(new_n557_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n588_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n625_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n590_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n591_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n616_), .B1(new_n662_), .B2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT98), .B1(new_n656_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n641_), .A2(new_n643_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n569_), .A2(new_n593_), .A3(new_n637_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n646_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n635_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n653_), .B1(new_n672_), .B2(new_n649_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n652_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n632_), .B1(new_n674_), .B2(new_n597_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT101), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT101), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n633_), .B1(new_n676_), .B2(new_n677_), .ZN(G1328gat));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n631_), .A2(new_n679_), .A3(new_n591_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT45), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n674_), .A2(new_n591_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n683_), .B2(G36gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT46), .ZN(G1329gat));
  INV_X1    g484(.A(G43gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n674_), .B2(new_n616_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n631_), .A2(new_n616_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1330gat));
  INV_X1    g490(.A(G50gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n631_), .A2(new_n692_), .A3(new_n527_), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT103), .B1(new_n674_), .B2(new_n527_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n695_), .B(new_n625_), .C1(new_n652_), .C2(new_n673_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT104), .B1(new_n697_), .B2(G50gat), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n699_));
  NOR4_X1   g498(.A1(new_n694_), .A2(new_n696_), .A3(new_n699_), .A4(new_n692_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n693_), .B1(new_n698_), .B2(new_n700_), .ZN(G1331gat));
  NOR2_X1   g500(.A1(new_n328_), .A2(new_n353_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n628_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n300_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n597_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n603_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n597_), .A2(G57gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1332gat));
  INV_X1    g509(.A(G64gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n704_), .A2(new_n711_), .A3(new_n591_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n708_), .A2(new_n591_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(G64gat), .ZN(new_n715_));
  AOI211_X1 g514(.A(KEYINPUT48), .B(new_n711_), .C1(new_n708_), .C2(new_n591_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT106), .ZN(G1333gat));
  AOI21_X1  g517(.A(new_n406_), .B1(new_n708_), .B2(new_n616_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT49), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n704_), .A2(new_n406_), .A3(new_n616_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1334gat));
  INV_X1    g521(.A(G78gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n708_), .B2(new_n527_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n704_), .A2(new_n723_), .A3(new_n527_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1335gat));
  INV_X1    g527(.A(new_n602_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n702_), .A2(new_n233_), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n729_), .B(new_n730_), .C1(new_n593_), .C2(new_n569_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n597_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n672_), .A2(new_n730_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n482_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(G1336gat));
  AOI21_X1  g534(.A(G92gat), .B1(new_n731_), .B2(new_n591_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n591_), .A2(G92gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n733_), .B2(new_n737_), .ZN(G1337gat));
  INV_X1    g537(.A(G99gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n733_), .B2(new_n616_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n731_), .A2(new_n269_), .A3(new_n616_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n742_));
  OAI22_X1  g541(.A1(new_n740_), .A2(new_n741_), .B1(new_n742_), .B2(KEYINPUT51), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(KEYINPUT51), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(G1338gat));
  NAND3_X1  g544(.A1(new_n731_), .A2(new_n270_), .A3(new_n527_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n270_), .B1(new_n733_), .B2(new_n527_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n747_), .A2(new_n748_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g551(.A1(new_n567_), .A2(new_n570_), .A3(new_n482_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n634_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n309_), .A2(KEYINPUT111), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT111), .B1(new_n309_), .B2(new_n756_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT12), .ZN(new_n759_));
  AOI211_X1 g558(.A(new_n759_), .B(new_n219_), .C1(new_n264_), .C2(new_n273_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n308_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n311_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n302_), .A2(KEYINPUT55), .A3(new_n303_), .A4(new_n308_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n757_), .A2(new_n758_), .A3(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n318_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n309_), .A2(new_n756_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n309_), .A2(KEYINPUT111), .A3(new_n756_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n769_), .A2(new_n763_), .A3(new_n762_), .A4(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n319_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n333_), .B1(new_n330_), .B2(new_n339_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n331_), .B(KEYINPUT113), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n344_), .B(new_n774_), .C1(new_n775_), .C2(new_n333_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n352_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n766_), .A2(new_n773_), .A3(new_n777_), .A4(new_n321_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n778_), .A2(KEYINPUT114), .A3(KEYINPUT58), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT58), .B1(new_n778_), .B2(KEYINPUT114), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n755_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT112), .B(KEYINPUT56), .C1(new_n765_), .C2(new_n318_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n320_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n771_), .B2(new_n319_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n784_), .B(new_n785_), .C1(new_n787_), .C2(KEYINPUT56), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n777_), .A2(new_n323_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT57), .B1(new_n790_), .B2(new_n729_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n792_), .B(new_n602_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT115), .B(new_n755_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n783_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n233_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n299_), .A2(new_n328_), .A3(new_n354_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT54), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT109), .B(KEYINPUT110), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n299_), .A2(new_n801_), .A3(new_n328_), .A4(new_n354_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n799_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n800_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n754_), .B1(new_n797_), .B2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(G113gat), .B1(new_n806_), .B2(new_n353_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n806_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n602_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT57), .ZN(new_n810_));
  INV_X1    g609(.A(new_n781_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n233_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n805_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n754_), .A2(KEYINPUT59), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n808_), .A2(KEYINPUT59), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n354_), .A2(new_n420_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n807_), .B1(new_n815_), .B2(new_n816_), .ZN(G1340gat));
  NAND2_X1  g616(.A1(new_n813_), .A2(new_n814_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n818_), .B(new_n329_), .C1(new_n806_), .C2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(G120gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n418_), .B1(new_n328_), .B2(KEYINPUT60), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n806_), .B(new_n822_), .C1(KEYINPUT60), .C2(new_n418_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT116), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n821_), .A2(new_n823_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n806_), .B2(new_n629_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n629_), .A2(G127gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT117), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n815_), .B2(new_n831_), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(new_n806_), .B2(new_n602_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n755_), .A2(G134gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n815_), .B2(new_n834_), .ZN(G1343gat));
  NAND3_X1  g634(.A1(new_n664_), .A2(new_n597_), .A3(new_n527_), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n616_), .B(new_n836_), .C1(new_n797_), .C2(new_n805_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n353_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT118), .B(G141gat), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(G1344gat));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n329_), .ZN(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT119), .B(G148gat), .Z(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1345gat));
  NAND2_X1  g642(.A1(new_n837_), .A2(new_n629_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G155gat), .ZN(new_n845_));
  INV_X1    g644(.A(G155gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n837_), .A2(new_n846_), .A3(new_n629_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n845_), .A2(new_n849_), .A3(new_n847_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1346gat));
  AOI21_X1  g652(.A(G162gat), .B1(new_n837_), .B2(new_n602_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n668_), .A2(G162gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n837_), .B2(new_n855_), .ZN(G1347gat));
  NAND2_X1  g655(.A1(new_n485_), .A2(new_n591_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT121), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n813_), .A2(new_n625_), .A3(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n354_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n356_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n860_), .A2(new_n354_), .A3(new_n538_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT62), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(KEYINPUT62), .B2(new_n862_), .ZN(G1348gat));
  AOI21_X1  g664(.A(new_n527_), .B1(new_n797_), .B2(new_n805_), .ZN(new_n866_));
  AND4_X1   g665(.A1(G176gat), .A2(new_n866_), .A3(new_n329_), .A4(new_n859_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n361_), .B1(new_n860_), .B2(new_n328_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n868_), .A2(KEYINPUT122), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(KEYINPUT122), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n869_), .B2(new_n870_), .ZN(G1349gat));
  NOR3_X1   g670(.A1(new_n860_), .A2(new_n392_), .A3(new_n233_), .ZN(new_n872_));
  INV_X1    g671(.A(G183gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n866_), .A2(new_n629_), .A3(new_n859_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(G1350gat));
  NAND2_X1  g674(.A1(new_n602_), .A2(new_n389_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n860_), .A2(new_n876_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n813_), .A2(new_n625_), .A3(new_n755_), .A4(new_n859_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n878_), .A2(new_n879_), .A3(G190gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n878_), .B2(G190gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n877_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n877_), .B(KEYINPUT124), .C1(new_n880_), .C2(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1351gat));
  AOI211_X1 g685(.A(new_n590_), .B(new_n616_), .C1(new_n797_), .C2(new_n805_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n887_), .A2(new_n591_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n353_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G197gat), .ZN(new_n890_));
  INV_X1    g689(.A(G197gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n888_), .A2(new_n891_), .A3(new_n353_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1352gat));
  NAND2_X1  g692(.A1(new_n888_), .A2(new_n329_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT125), .B(G204gat), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n888_), .A2(new_n329_), .A3(new_n895_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1353gat));
  NAND3_X1  g698(.A1(new_n887_), .A2(new_n591_), .A3(new_n629_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n901_), .ZN(G1354gat));
  AOI21_X1  g703(.A(new_n616_), .B1(new_n797_), .B2(new_n805_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n905_), .A2(new_n663_), .A3(new_n591_), .A4(new_n602_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n887_), .A2(KEYINPUT126), .A3(new_n591_), .A4(new_n602_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT127), .B(G218gat), .Z(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n908_), .A2(new_n909_), .A3(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n888_), .A2(new_n755_), .A3(new_n910_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1355gat));
endmodule


