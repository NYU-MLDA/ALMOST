//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n943_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n968_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n981_, new_n982_, new_n983_, new_n984_, new_n986_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n994_,
    new_n995_, new_n996_;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G127gat), .B(G134gat), .Z(new_n205_));
  XOR2_X1   g004(.A(G113gat), .B(G120gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR3_X1   g012(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT86), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n213_), .B1(new_n216_), .B2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n217_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n211_), .B1(KEYINPUT1), .B2(new_n209_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n208_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n214_), .A2(new_n215_), .ZN(new_n231_));
  NOR4_X1   g030(.A1(KEYINPUT86), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n222_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n229_), .B1(new_n233_), .B2(new_n212_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n207_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n235_), .A3(KEYINPUT4), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n234_), .A2(new_n207_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT96), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT96), .ZN(new_n240_));
  NOR4_X1   g039(.A1(new_n234_), .A2(new_n207_), .A3(new_n240_), .A4(KEYINPUT4), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n204_), .B(new_n236_), .C1(new_n239_), .C2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n230_), .A2(new_n235_), .A3(new_n203_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G1gat), .B(G29gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G85gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT0), .B(G57gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT100), .ZN(new_n250_));
  INV_X1    g049(.A(new_n248_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n242_), .A2(new_n243_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n249_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n244_), .A2(KEYINPUT100), .A3(new_n248_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G78gat), .B(G106gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n233_), .A2(new_n212_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n229_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT89), .ZN(new_n263_));
  INV_X1    g062(.A(G204gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(G197gat), .ZN(new_n265_));
  INV_X1    g064(.A(G197gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(G197gat), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n265_), .A2(new_n267_), .A3(new_n268_), .A4(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n264_), .A2(G197gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT21), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT90), .ZN(new_n275_));
  INV_X1    g074(.A(G218gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G211gat), .ZN(new_n277_));
  INV_X1    g076(.A(G211gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G218gat), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n277_), .A2(new_n279_), .A3(KEYINPUT90), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n270_), .B(new_n273_), .C1(new_n275_), .C2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n279_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT90), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n274_), .A2(KEYINPUT90), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n265_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(KEYINPUT21), .A4(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT88), .B1(new_n262_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G228gat), .A2(G233gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT88), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n293_), .B(new_n288_), .C1(new_n234_), .C2(new_n259_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n290_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n292_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n258_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT91), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n234_), .A2(new_n259_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G22gat), .B(G50gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n300_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n294_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT29), .B1(new_n223_), .B2(new_n229_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n293_), .B1(new_n306_), .B2(new_n288_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n291_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n290_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n257_), .A3(new_n309_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n299_), .A2(new_n304_), .B1(new_n297_), .B2(new_n310_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n297_), .A2(KEYINPUT91), .A3(new_n310_), .A4(new_n304_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G71gat), .B(G99gat), .ZN(new_n314_));
  INV_X1    g113(.A(G43gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT30), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(G183gat), .A3(G190gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n319_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT81), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n324_), .A2(new_n325_), .A3(KEYINPUT23), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n324_), .B2(KEYINPUT23), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n322_), .B(new_n323_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT26), .B(G190gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT79), .B1(new_n330_), .B2(G183gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT25), .B(G183gat), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n329_), .B(new_n331_), .C1(new_n332_), .C2(KEYINPUT79), .ZN(new_n333_));
  OR3_X1    g132(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT80), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G169gat), .A3(G176gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n338_), .A3(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n328_), .A2(new_n333_), .A3(new_n334_), .A4(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT83), .B(G15gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G169gat), .ZN(new_n347_));
  INV_X1    g146(.A(G176gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n338_), .A2(new_n340_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n320_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n319_), .B1(G183gat), .B2(G190gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n349_), .B(new_n350_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n342_), .A2(new_n346_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n346_), .B1(new_n342_), .B2(new_n355_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n318_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n342_), .A2(new_n355_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n345_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n316_), .B(KEYINPUT30), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(new_n356_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n359_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n359_), .B2(new_n363_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n207_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n359_), .A2(new_n363_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n364_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n359_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n208_), .A3(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n368_), .A2(new_n372_), .A3(KEYINPUT85), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT85), .B1(new_n368_), .B2(new_n372_), .ZN(new_n374_));
  OAI22_X1  g173(.A1(new_n311_), .A2(new_n313_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n257_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n304_), .B1(new_n376_), .B2(KEYINPUT91), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n297_), .A2(new_n310_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n368_), .A2(new_n372_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n312_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n256_), .B1(new_n375_), .B2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT18), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n328_), .B1(G183gat), .B2(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n349_), .A2(new_n350_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT94), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT94), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n351_), .A2(new_n352_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n332_), .A2(new_n329_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n336_), .A2(new_n337_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n397_), .A2(new_n334_), .A3(new_n398_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n390_), .B1(new_n401_), .B2(new_n288_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n360_), .A2(new_n288_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT20), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT95), .ZN(new_n406_));
  AND4_X1   g205(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .A4(new_n334_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT94), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT94), .B1(new_n349_), .B2(new_n350_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n407_), .B1(new_n410_), .B2(new_n391_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n406_), .B1(new_n411_), .B2(new_n289_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT20), .B1(new_n360_), .B2(new_n288_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT93), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n401_), .A2(KEYINPUT95), .A3(new_n288_), .ZN(new_n416_));
  OAI211_X1 g215(.A(KEYINPUT93), .B(KEYINPUT20), .C1(new_n360_), .C2(new_n288_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n412_), .A2(new_n415_), .A3(new_n416_), .A4(new_n417_), .ZN(new_n418_));
  AOI211_X1 g217(.A(new_n386_), .B(new_n405_), .C1(new_n389_), .C2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT101), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n418_), .A2(new_n389_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n411_), .A2(KEYINPUT99), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT99), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n401_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n424_), .A3(new_n289_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n404_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n390_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n421_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n386_), .ZN(new_n429_));
  OAI22_X1  g228(.A1(new_n419_), .A2(new_n420_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n405_), .B1(new_n418_), .B2(new_n389_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n429_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(KEYINPUT101), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT27), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n431_), .A2(new_n429_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT27), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n432_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT97), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n242_), .A2(new_n243_), .A3(new_n251_), .A4(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n203_), .B(new_n236_), .C1(new_n239_), .C2(new_n241_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n230_), .A2(new_n235_), .A3(new_n204_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n248_), .A3(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n252_), .A2(KEYINPUT97), .A3(new_n439_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n435_), .A2(new_n445_), .A3(new_n432_), .A4(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT98), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n429_), .A2(KEYINPUT32), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n431_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n431_), .B2(new_n449_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(KEYINPUT32), .B(new_n429_), .C1(new_n421_), .C2(new_n427_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n253_), .A2(new_n453_), .A3(new_n254_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n447_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n373_), .A2(new_n374_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n379_), .A2(new_n312_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n382_), .A2(new_n438_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G15gat), .B(G22gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G1gat), .A2(G8gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT14), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(G1gat), .A2(G8gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n461_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n460_), .A2(new_n461_), .A3(new_n464_), .A4(new_n462_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G29gat), .B(G36gat), .Z(new_n472_));
  XOR2_X1   g271(.A(G43gat), .B(G50gat), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n468_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n471_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT15), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n474_), .A2(KEYINPUT15), .A3(new_n471_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n468_), .A3(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n479_), .A3(new_n477_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n481_), .A2(new_n486_), .A3(KEYINPUT77), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT77), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n478_), .A2(new_n488_), .A3(new_n480_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G113gat), .B(G141gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G169gat), .B(G197gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(KEYINPUT78), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n487_), .B(new_n489_), .C1(KEYINPUT78), .C2(new_n494_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n202_), .B1(new_n459_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n455_), .A2(new_n458_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n368_), .A2(new_n372_), .A3(KEYINPUT85), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n380_), .A2(new_n502_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n501_), .A2(new_n503_), .B1(new_n379_), .B2(new_n312_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n379_), .A2(new_n312_), .A3(new_n380_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n255_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n435_), .A2(new_n436_), .A3(new_n432_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n419_), .A2(new_n420_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n432_), .A2(KEYINPUT101), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n508_), .B(new_n509_), .C1(new_n429_), .C2(new_n428_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n507_), .B1(new_n510_), .B2(KEYINPUT27), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n500_), .B1(new_n506_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n498_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(KEYINPUT102), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n499_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G190gat), .B(G218gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G134gat), .B(G162gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT36), .Z(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT10), .B(G99gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT64), .B(G106gat), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT6), .ZN(new_n524_));
  INV_X1    g323(.A(G85gat), .ZN(new_n525_));
  INV_X1    g324(.A(G92gat), .ZN(new_n526_));
  OR3_X1    g325(.A1(new_n525_), .A2(new_n526_), .A3(KEYINPUT9), .ZN(new_n527_));
  XOR2_X1   g326(.A(G85gat), .B(G92gat), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT9), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n522_), .A2(new_n524_), .A3(new_n527_), .A4(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT8), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT66), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT6), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT66), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n523_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(KEYINPUT65), .A2(G99gat), .ZN(new_n537_));
  INV_X1    g336(.A(G106gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT7), .ZN(new_n540_));
  NOR3_X1   g339(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT7), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n534_), .A2(KEYINPUT66), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n532_), .A2(KEYINPUT6), .ZN(new_n545_));
  AND2_X1   g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n536_), .A2(new_n540_), .A3(new_n543_), .A4(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n531_), .B1(new_n548_), .B2(new_n528_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n528_), .A2(new_n531_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n541_), .B(KEYINPUT7), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n551_), .B2(new_n524_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n530_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT67), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(KEYINPUT67), .B(new_n530_), .C1(new_n549_), .C2(new_n552_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n476_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT35), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n483_), .A2(new_n484_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n553_), .A2(new_n564_), .B1(new_n561_), .B2(new_n560_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n557_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n563_), .B1(new_n557_), .B2(new_n565_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n519_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n518_), .A2(KEYINPUT36), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n566_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n569_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT72), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT72), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n569_), .A2(new_n572_), .A3(new_n576_), .A4(new_n573_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n569_), .A2(KEYINPUT71), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n572_), .B1(new_n569_), .B2(KEYINPUT71), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT37), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n468_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G71gat), .B(G78gat), .Z(new_n586_));
  INV_X1    g385(.A(G64gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(G57gat), .ZN(new_n588_));
  INV_X1    g387(.A(G57gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(G64gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n590_), .A3(KEYINPUT11), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n588_), .A2(new_n590_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(KEYINPUT11), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n586_), .A2(new_n591_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n592_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n466_), .A2(new_n467_), .A3(new_n583_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n585_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n592_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n593_), .A2(KEYINPUT11), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n600_), .B1(new_n601_), .B2(new_n595_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n466_), .A2(new_n467_), .A3(new_n583_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n583_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n602_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT73), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n599_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n608_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n609_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n608_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n611_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n607_), .A2(KEYINPUT17), .A3(new_n612_), .A4(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n606_), .B1(new_n599_), .B2(new_n605_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT17), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n617_), .A2(new_n618_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n610_), .A2(new_n611_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n623_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n619_), .A2(new_n612_), .A3(KEYINPUT17), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT75), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n599_), .A2(new_n605_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n599_), .B2(new_n605_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n628_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT76), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n628_), .B(KEYINPUT76), .C1(new_n630_), .C2(new_n631_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n622_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n582_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(G230gat), .ZN(new_n638_));
  INV_X1    g437(.A(G233gat), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n555_), .A2(new_n602_), .A3(new_n556_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n602_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n553_), .A2(KEYINPUT12), .A3(new_n597_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n642_), .B2(KEYINPUT12), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n555_), .A2(new_n602_), .A3(new_n556_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n640_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n643_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(G120gat), .B(G148gat), .Z(new_n650_));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT68), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT70), .Z(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n649_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n656_), .B(new_n643_), .C1(new_n645_), .C2(new_n648_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT13), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(KEYINPUT13), .A3(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n637_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n255_), .A2(G1gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n515_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT103), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(KEYINPUT103), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT38), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n569_), .A2(new_n572_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n459_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n636_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n664_), .A2(new_n498_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT104), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n675_), .A2(new_n680_), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n256_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G1gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n668_), .A2(KEYINPUT38), .A3(new_n669_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n672_), .A2(new_n684_), .A3(new_n685_), .ZN(G1324gat));
  AND2_X1   g485(.A1(new_n515_), .A2(new_n665_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n438_), .A2(G8gat), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT39), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n512_), .A2(new_n511_), .A3(new_n673_), .A4(new_n677_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT105), .B1(new_n690_), .B2(G8gat), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n687_), .A2(new_n688_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n689_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n690_), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1325gat));
  INV_X1    g497(.A(G15gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n687_), .A2(new_n699_), .A3(new_n456_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n682_), .B2(new_n456_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT41), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT41), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n702_), .B2(new_n703_), .ZN(G1326gat));
  INV_X1    g503(.A(G22gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n687_), .A2(new_n705_), .A3(new_n457_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n682_), .A2(new_n457_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(G22gat), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT42), .B(new_n705_), .C1(new_n682_), .C2(new_n457_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(G1327gat));
  NAND2_X1  g510(.A1(new_n674_), .A2(new_n676_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n664_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n499_), .B2(new_n514_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G29gat), .B1(new_n715_), .B2(new_n256_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n459_), .B2(new_n582_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n718_));
  INV_X1    g517(.A(new_n582_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n512_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n664_), .A2(new_n498_), .A3(new_n636_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT44), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724_));
  INV_X1    g523(.A(new_n722_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n724_), .B(new_n725_), .C1(new_n717_), .C2(new_n720_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n723_), .A2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n256_), .A2(G29gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n716_), .B1(new_n727_), .B2(new_n728_), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n727_), .B2(new_n511_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n438_), .A2(KEYINPUT107), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n438_), .A2(KEYINPUT107), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(G36gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n515_), .A2(new_n713_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT45), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n715_), .A2(new_n739_), .A3(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n730_), .B1(new_n732_), .B2(new_n742_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n723_), .A2(new_n726_), .A3(new_n438_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n741_), .B(KEYINPUT46), .C1(new_n744_), .C2(new_n731_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1329gat));
  INV_X1    g545(.A(new_n380_), .ZN(new_n747_));
  NOR4_X1   g546(.A1(new_n723_), .A2(new_n726_), .A3(new_n315_), .A4(new_n747_), .ZN(new_n748_));
  XOR2_X1   g547(.A(KEYINPUT108), .B(G43gat), .Z(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n715_), .B2(new_n456_), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT47), .B1(new_n748_), .B2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n727_), .A2(G43gat), .A3(new_n380_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n750_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n751_), .A2(new_n755_), .ZN(G1330gat));
  AOI21_X1  g555(.A(G50gat), .B1(new_n715_), .B2(new_n457_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n457_), .A2(G50gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n727_), .B2(new_n758_), .ZN(G1331gat));
  NOR2_X1   g558(.A1(new_n459_), .A2(new_n513_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n582_), .A2(new_n664_), .A3(new_n636_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G57gat), .B1(new_n764_), .B2(new_n256_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n589_), .B1(new_n256_), .B2(KEYINPUT110), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n675_), .A2(new_n498_), .A3(new_n664_), .A4(new_n636_), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n766_), .B(new_n767_), .C1(KEYINPUT110), .C2(new_n589_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n765_), .A2(new_n768_), .ZN(G1332gat));
  OAI21_X1  g568(.A(G64gat), .B1(new_n767_), .B2(new_n735_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT48), .ZN(new_n771_));
  INV_X1    g570(.A(new_n735_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n764_), .A2(new_n587_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1333gat));
  INV_X1    g573(.A(new_n456_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G71gat), .B1(new_n767_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT49), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n775_), .A2(G71gat), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT111), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n764_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1334gat));
  INV_X1    g580(.A(new_n457_), .ZN(new_n782_));
  OAI21_X1  g581(.A(G78gat), .B1(new_n767_), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT50), .ZN(new_n784_));
  INV_X1    g583(.A(G78gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n764_), .A2(new_n785_), .A3(new_n457_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1335gat));
  INV_X1    g586(.A(new_n664_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n788_), .A2(new_n513_), .A3(new_n636_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n721_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n255_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n788_), .A2(new_n712_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n760_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n525_), .A3(new_n256_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(new_n795_), .ZN(G1336gat));
  OAI21_X1  g595(.A(new_n526_), .B1(new_n793_), .B2(new_n438_), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT112), .Z(new_n798_));
  NOR3_X1   g597(.A1(new_n790_), .A2(new_n526_), .A3(new_n735_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n790_), .B2(new_n775_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n747_), .A2(new_n520_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n793_), .B2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g603(.A1(new_n793_), .A2(new_n782_), .A3(new_n521_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n721_), .A2(new_n457_), .A3(new_n789_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n538_), .B1(new_n807_), .B2(KEYINPUT52), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(KEYINPUT52), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n806_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n805_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT53), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n814_), .B(new_n805_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(G1339gat));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n634_), .A2(new_n635_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n622_), .ZN(new_n822_));
  AND4_X1   g621(.A1(KEYINPUT114), .A2(new_n821_), .A3(new_n498_), .A4(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT114), .B1(new_n636_), .B2(new_n498_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n826_), .A2(KEYINPUT115), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n825_), .A2(new_n662_), .A3(new_n828_), .A4(new_n663_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n582_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n820_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n826_), .A2(KEYINPUT115), .ZN(new_n832_));
  INV_X1    g631(.A(new_n820_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n582_), .A3(new_n833_), .A4(new_n829_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n819_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n490_), .A2(new_n494_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n494_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT118), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n485_), .A2(new_n477_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n840_), .A2(KEYINPUT119), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n479_), .B1(new_n840_), .B2(KEYINPUT119), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n837_), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n659_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n646_), .A2(new_n647_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n524_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n540_), .A2(new_n543_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n531_), .B(new_n528_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n528_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n546_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n851_), .B1(new_n854_), .B2(new_n551_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n850_), .B1(new_n855_), .B2(new_n531_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT67), .B1(new_n856_), .B2(new_n530_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n556_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n597_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT12), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n847_), .A2(new_n861_), .A3(new_n644_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n656_), .B1(new_n862_), .B2(new_n643_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n845_), .B1(new_n846_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n844_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT120), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n870_));
  INV_X1    g669(.A(new_n654_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n646_), .B(new_n644_), .C1(new_n642_), .C2(KEYINPUT12), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n862_), .A2(new_n872_), .B1(new_n640_), .B2(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n847_), .A2(new_n861_), .A3(KEYINPUT55), .A4(new_n644_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n871_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n870_), .B1(new_n876_), .B2(KEYINPUT117), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n643_), .B(new_n871_), .C1(new_n645_), .C2(new_n648_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n513_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n872_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n873_), .A2(new_n640_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n875_), .A3(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT117), .B1(new_n882_), .B2(new_n654_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n879_), .B1(new_n883_), .B2(KEYINPUT56), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n869_), .B1(new_n877_), .B2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n836_), .B1(new_n885_), .B2(new_n674_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n877_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n867_), .B(new_n865_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n674_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT57), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n882_), .A2(new_n654_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT56), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n882_), .A2(new_n870_), .A3(new_n654_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n845_), .A2(new_n878_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n892_), .A2(KEYINPUT58), .A3(new_n893_), .A4(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n893_), .A2(new_n894_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n898_), .A2(KEYINPUT121), .A3(KEYINPUT58), .A4(new_n892_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n893_), .A2(new_n894_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n870_), .B1(new_n882_), .B2(new_n654_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n897_), .A2(new_n899_), .A3(new_n719_), .A4(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n886_), .A2(new_n890_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n835_), .B1(new_n905_), .B2(new_n676_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n511_), .A2(new_n255_), .A3(new_n381_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT59), .B1(new_n906_), .B2(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n904_), .B1(KEYINPUT57), .B2(new_n889_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n885_), .A2(new_n836_), .A3(new_n674_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n676_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n835_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n908_), .A2(KEYINPUT122), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n908_), .A2(KEYINPUT122), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n915_), .A2(new_n916_), .A3(KEYINPUT59), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n914_), .A2(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n909_), .A2(new_n513_), .A3(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G113gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n914_), .A2(new_n907_), .ZN(new_n921_));
  OR3_X1    g720(.A1(new_n921_), .A2(G113gat), .A3(new_n498_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n922_), .ZN(G1340gat));
  NAND3_X1  g722(.A1(new_n909_), .A2(new_n664_), .A3(new_n918_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G120gat), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n906_), .A2(new_n908_), .ZN(new_n926_));
  INV_X1    g725(.A(G120gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n788_), .B2(KEYINPUT60), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n926_), .B(new_n928_), .C1(KEYINPUT60), .C2(new_n927_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n929_), .ZN(G1341gat));
  NAND3_X1  g729(.A1(new_n909_), .A2(new_n636_), .A3(new_n918_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(G127gat), .ZN(new_n932_));
  OR3_X1    g731(.A1(new_n921_), .A2(G127gat), .A3(new_n676_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1342gat));
  AOI21_X1  g733(.A(G134gat), .B1(new_n926_), .B2(new_n674_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n909_), .A2(new_n918_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n719_), .A2(G134gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT123), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n935_), .B1(new_n936_), .B2(new_n938_), .ZN(G1343gat));
  NOR3_X1   g738(.A1(new_n772_), .A2(new_n255_), .A3(new_n375_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n914_), .A2(new_n513_), .A3(new_n940_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g741(.A1(new_n914_), .A2(new_n664_), .A3(new_n940_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g743(.A1(new_n914_), .A2(new_n636_), .A3(new_n940_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(KEYINPUT61), .B(G155gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(G1346gat));
  INV_X1    g746(.A(G162gat), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n914_), .A2(new_n948_), .A3(new_n674_), .A4(new_n940_), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n914_), .A2(new_n719_), .A3(new_n940_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n948_), .ZN(G1347gat));
  AND2_X1   g750(.A1(new_n513_), .A2(new_n347_), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n772_), .A2(new_n255_), .A3(new_n782_), .A4(new_n456_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(KEYINPUT124), .B1(new_n914_), .B2(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n906_), .A2(new_n956_), .A3(new_n953_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n952_), .B1(new_n955_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(G169gat), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n953_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n960_));
  AOI211_X1 g759(.A(KEYINPUT62), .B(new_n959_), .C1(new_n960_), .C2(new_n513_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n914_), .A2(new_n513_), .A3(new_n954_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n962_), .B1(new_n963_), .B2(G169gat), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n958_), .B1(new_n961_), .B2(new_n964_), .ZN(G1348gat));
  OAI211_X1 g764(.A(new_n348_), .B(new_n664_), .C1(new_n955_), .C2(new_n957_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n960_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G176gat), .B1(new_n967_), .B2(new_n788_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n966_), .A2(new_n968_), .ZN(G1349gat));
  AOI21_X1  g768(.A(G183gat), .B1(new_n960_), .B2(new_n636_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n960_), .A2(KEYINPUT124), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n956_), .B1(new_n906_), .B2(new_n953_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n971_), .A2(new_n972_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n676_), .A2(new_n332_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n970_), .B1(new_n973_), .B2(new_n974_), .ZN(G1350gat));
  AND2_X1   g774(.A1(new_n674_), .A2(new_n329_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n976_), .B1(new_n955_), .B2(new_n957_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n582_), .B1(new_n971_), .B2(new_n972_), .ZN(new_n978_));
  INV_X1    g777(.A(G190gat), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n977_), .B1(new_n978_), .B2(new_n979_), .ZN(G1351gat));
  NOR3_X1   g779(.A1(new_n735_), .A2(new_n256_), .A3(new_n375_), .ZN(new_n981_));
  AND2_X1   g780(.A1(new_n914_), .A2(new_n981_), .ZN(new_n982_));
  AOI21_X1  g781(.A(G197gat), .B1(new_n982_), .B2(new_n513_), .ZN(new_n983_));
  AND4_X1   g782(.A1(G197gat), .A2(new_n914_), .A3(new_n513_), .A4(new_n981_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n983_), .A2(new_n984_), .ZN(G1352gat));
  NAND3_X1  g784(.A1(new_n914_), .A2(new_n664_), .A3(new_n981_), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n986_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g786(.A(new_n676_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n988_));
  XOR2_X1   g787(.A(new_n988_), .B(KEYINPUT125), .Z(new_n989_));
  NAND3_X1  g788(.A1(new_n914_), .A2(new_n981_), .A3(new_n989_), .ZN(new_n990_));
  NOR2_X1   g789(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n991_));
  XOR2_X1   g790(.A(new_n991_), .B(KEYINPUT126), .Z(new_n992_));
  XNOR2_X1  g791(.A(new_n990_), .B(new_n992_), .ZN(G1354gat));
  NAND2_X1  g792(.A1(new_n982_), .A2(new_n674_), .ZN(new_n994_));
  XNOR2_X1  g793(.A(KEYINPUT127), .B(G218gat), .ZN(new_n995_));
  NOR2_X1   g794(.A1(new_n582_), .A2(new_n995_), .ZN(new_n996_));
  AOI22_X1  g795(.A1(new_n994_), .A2(new_n995_), .B1(new_n982_), .B2(new_n996_), .ZN(G1355gat));
endmodule


