//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n553_, new_n554_, new_n555_, new_n556_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT75), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT74), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n213_), .B(KEYINPUT23), .Z(new_n214_));
  NOR2_X1   g013(.A1(new_n209_), .A2(KEYINPUT24), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(G190gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT26), .B1(new_n218_), .B2(KEYINPUT73), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(KEYINPUT26), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n217_), .B(new_n219_), .C1(new_n220_), .C2(KEYINPUT73), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n212_), .A2(new_n216_), .A3(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT22), .B(G169gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n208_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n224_), .B(new_n210_), .C1(new_n214_), .C2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n206_), .B(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G227gat), .A2(G233gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G71gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(G15gat), .B(G43gat), .Z(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT30), .B(G99gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n228_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237_));
  AND2_X1   g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT77), .B1(KEYINPUT76), .B2(KEYINPUT3), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G141gat), .A2(G148gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n241_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(new_n242_), .B2(new_n241_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n246_), .B(KEYINPUT2), .Z(new_n247_));
  OAI21_X1  g046(.A(new_n240_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n239_), .B1(new_n238_), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n249_), .B2(new_n238_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n242_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(new_n252_), .A3(new_n246_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n237_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G211gat), .B(G218gat), .ZN(new_n255_));
  INV_X1    g054(.A(G197gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT79), .B1(new_n256_), .B2(G204gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(KEYINPUT21), .A3(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G197gat), .B(G204gat), .Z(new_n259_));
  OR2_X1    g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n258_), .B(new_n259_), .C1(KEYINPUT21), .C2(new_n255_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(G228gat), .B(G233gat), .C1(new_n254_), .C2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G228gat), .A2(G233gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n261_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n248_), .A2(new_n253_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n264_), .B(new_n265_), .C1(new_n266_), .C2(new_n237_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G78gat), .B(G106gat), .Z(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n248_), .A2(new_n253_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(KEYINPUT29), .ZN(new_n273_));
  XOR2_X1   g072(.A(G22gat), .B(G50gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT78), .B(KEYINPUT28), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n273_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n263_), .A2(new_n267_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n268_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n269_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n278_), .A2(new_n282_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n204_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n272_), .A2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(KEYINPUT4), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n248_), .A2(new_n253_), .A3(new_n204_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n266_), .A2(KEYINPUT86), .A3(new_n204_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n289_), .B1(new_n294_), .B2(KEYINPUT4), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(KEYINPUT87), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n297_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(KEYINPUT88), .B(KEYINPUT0), .Z(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G29gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G57gat), .B(G85gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n306_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n298_), .A2(new_n308_), .A3(new_n300_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n227_), .A2(new_n265_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT82), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n227_), .A2(KEYINPUT82), .A3(new_n265_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT26), .B(G190gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n217_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n216_), .A2(new_n211_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n226_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(new_n265_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(KEYINPUT83), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n320_), .B2(KEYINPUT83), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n315_), .A2(new_n321_), .A3(new_n324_), .A4(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT85), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT32), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n325_), .B1(new_n319_), .B2(new_n265_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n265_), .B2(new_n227_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n324_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n327_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n336_), .A2(new_n337_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n320_), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n342_));
  NAND3_X1  g141(.A1(new_n315_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n340_), .B1(new_n343_), .B2(new_n337_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(new_n334_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n310_), .A2(new_n339_), .A3(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n327_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n333_), .B1(new_n327_), .B2(new_n338_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n295_), .A2(new_n299_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n294_), .A2(new_n297_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n306_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT33), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n309_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n298_), .A2(KEYINPUT33), .A3(new_n308_), .A4(new_n300_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n349_), .A2(new_n352_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n286_), .B1(new_n346_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n327_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(KEYINPUT27), .C1(new_n344_), .C2(new_n333_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n362_), .A2(new_n310_), .A3(new_n285_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n236_), .B1(new_n357_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n362_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT90), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n307_), .A2(new_n309_), .A3(new_n235_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n365_), .A2(new_n366_), .A3(new_n285_), .A4(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n359_), .A2(new_n285_), .A3(new_n361_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT90), .B1(new_n370_), .B2(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n364_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G71gat), .B(G78gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G57gat), .B(G64gat), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(KEYINPUT11), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(KEYINPUT11), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n374_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n377_), .A2(new_n374_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT12), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT65), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT65), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT6), .ZN(new_n387_));
  AND2_X1   g186(.A1(G99gat), .A2(G106gat), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n385_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n388_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT7), .ZN(new_n391_));
  INV_X1    g190(.A(G99gat), .ZN(new_n392_));
  INV_X1    g191(.A(G106gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n389_), .A2(new_n390_), .A3(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G85gat), .B(G92gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT67), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT8), .B1(new_n397_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT8), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n385_), .A2(new_n387_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n388_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n385_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n403_), .B(new_n400_), .C1(new_n408_), .C2(new_n396_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n402_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n411_), .A2(G99gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n392_), .A2(KEYINPUT10), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n393_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  AND4_X1   g213(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n406_), .A2(new_n414_), .A3(new_n407_), .A4(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n418_));
  AOI211_X1 g217(.A(KEYINPUT64), .B(new_n418_), .C1(new_n398_), .C2(KEYINPUT9), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT66), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n389_), .A2(new_n390_), .ZN(new_n421_));
  AND2_X1   g220(.A1(G85gat), .A2(G92gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(G85gat), .A2(G92gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT9), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT64), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n424_), .B(new_n425_), .C1(KEYINPUT9), .C2(new_n422_), .ZN(new_n426_));
  XOR2_X1   g225(.A(KEYINPUT10), .B(G99gat), .Z(new_n427_));
  AOI21_X1  g226(.A(new_n415_), .B1(new_n427_), .B2(new_n393_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT66), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n421_), .A2(new_n426_), .A3(new_n428_), .A4(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n420_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT68), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n410_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n410_), .B2(new_n431_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n383_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n410_), .A2(new_n431_), .A3(new_n380_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT12), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n410_), .A2(new_n431_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n381_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G230gat), .A2(G233gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n435_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n436_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n441_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n446_));
  XNOR2_X1  g245(.A(G120gat), .B(G148gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G176gat), .B(G204gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n442_), .A2(new_n445_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT70), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT70), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n442_), .A2(new_n454_), .A3(new_n445_), .A4(new_n451_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n442_), .A2(new_n445_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n450_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(KEYINPUT13), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT13), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G29gat), .B(G36gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G43gat), .B(G50gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT72), .Z(new_n467_));
  XNOR2_X1  g266(.A(G15gat), .B(G22gat), .ZN(new_n468_));
  INV_X1    g267(.A(G1gat), .ZN(new_n469_));
  INV_X1    g268(.A(G8gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT14), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G1gat), .B(G8gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n467_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n476_));
  XNOR2_X1  g275(.A(new_n466_), .B(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n467_), .B(new_n474_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n479_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G113gat), .B(G141gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G169gat), .B(G197gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n463_), .A2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n373_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G231gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n474_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(new_n380_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G127gat), .B(G155gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G211gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT16), .B(G183gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n500_), .A2(KEYINPUT17), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n500_), .A2(KEYINPUT17), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n496_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n477_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n410_), .A2(new_n431_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT35), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G232gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT34), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n507_), .A2(new_n466_), .B1(new_n508_), .B2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n508_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n506_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n506_), .B2(new_n512_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G190gat), .B(G218gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G134gat), .B(G162gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(KEYINPUT36), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n520_), .B(KEYINPUT36), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT37), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n493_), .A2(new_n505_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(new_n469_), .A3(new_n310_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT38), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n460_), .A2(new_n462_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(new_n490_), .A3(new_n505_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n526_), .B(new_n373_), .C1(new_n533_), .C2(KEYINPUT91), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(KEYINPUT91), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT92), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n538_), .A2(new_n310_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n531_), .B1(new_n539_), .B2(new_n469_), .ZN(G1324gat));
  NOR3_X1   g339(.A1(new_n528_), .A2(G8gat), .A3(new_n365_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n537_), .B2(new_n365_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n535_), .A2(KEYINPUT93), .A3(new_n536_), .A4(new_n362_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(G8gat), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT39), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT39), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n543_), .A2(new_n547_), .A3(G8gat), .A4(new_n544_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n541_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT94), .B(KEYINPUT40), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n549_), .B(new_n551_), .ZN(G1325gat));
  INV_X1    g351(.A(G15gat), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n538_), .B2(new_n235_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT41), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n529_), .A2(new_n553_), .A3(new_n235_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(G1326gat));
  INV_X1    g356(.A(G22gat), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n538_), .B2(new_n286_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT42), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n286_), .A2(new_n558_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT95), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n528_), .B2(new_n563_), .ZN(G1327gat));
  INV_X1    g363(.A(G29gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n505_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n527_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT96), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT43), .B1(new_n527_), .B2(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n373_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n373_), .B2(new_n567_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n492_), .B(new_n566_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT44), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n527_), .B1(new_n364_), .B2(new_n372_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(new_n569_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(KEYINPUT44), .A3(new_n492_), .A4(new_n566_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n565_), .B1(new_n578_), .B2(new_n310_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n526_), .A2(new_n505_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT97), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n493_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n310_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n582_), .A2(G29gat), .A3(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n579_), .A2(new_n584_), .ZN(G1328gat));
  NAND3_X1  g384(.A1(new_n574_), .A2(new_n577_), .A3(new_n362_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n574_), .A2(new_n577_), .A3(KEYINPUT98), .A4(new_n362_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(G36gat), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n362_), .B(KEYINPUT99), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n582_), .A2(G36gat), .A3(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT100), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT45), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n593_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT45), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n590_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT46), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n590_), .A2(new_n595_), .A3(new_n599_), .A4(KEYINPUT46), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1329gat));
  NAND3_X1  g403(.A1(new_n578_), .A2(G43gat), .A3(new_n235_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n582_), .A2(new_n236_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(G43gat), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g407(.A1(new_n578_), .A2(new_n286_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(G50gat), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n285_), .A2(G50gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT101), .Z(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n582_), .B2(new_n612_), .ZN(G1331gat));
  AOI21_X1  g412(.A(new_n490_), .B1(new_n364_), .B2(new_n372_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n463_), .A2(new_n527_), .A3(new_n505_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n614_), .B1(KEYINPUT102), .B2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(KEYINPUT102), .B2(new_n615_), .ZN(new_n617_));
  AOI21_X1  g416(.A(G57gat), .B1(new_n617_), .B2(new_n310_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT103), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n614_), .A2(new_n463_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n505_), .A3(new_n526_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n310_), .A2(G57gat), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n619_), .B1(new_n622_), .B2(new_n623_), .ZN(G1332gat));
  OAI21_X1  g423(.A(G64gat), .B1(new_n621_), .B2(new_n592_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT48), .ZN(new_n626_));
  INV_X1    g425(.A(G64gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n617_), .A2(new_n627_), .A3(new_n591_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1333gat));
  INV_X1    g428(.A(G71gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n617_), .A2(new_n630_), .A3(new_n235_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n622_), .B2(new_n235_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT104), .B(KEYINPUT49), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n632_), .A2(new_n633_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n631_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT105), .ZN(G1334gat));
  OAI21_X1  g437(.A(G78gat), .B1(new_n621_), .B2(new_n285_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT106), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT50), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n641_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n285_), .A2(G78gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT107), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n617_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(new_n643_), .A3(new_n646_), .ZN(G1335gat));
  NAND2_X1  g446(.A1(new_n620_), .A2(new_n581_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n648_), .A2(G85gat), .A3(new_n583_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n532_), .A2(new_n490_), .A3(new_n505_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n576_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n310_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n649_), .B1(new_n652_), .B2(G85gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT108), .ZN(G1336gat));
  INV_X1    g453(.A(G92gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n655_), .B1(new_n648_), .B2(new_n365_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT109), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n592_), .A2(new_n655_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n651_), .B2(new_n658_), .ZN(G1337gat));
  INV_X1    g458(.A(KEYINPUT113), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT111), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n235_), .A2(new_n427_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n620_), .A2(new_n581_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n235_), .B(new_n650_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT110), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n665_), .A2(new_n666_), .A3(G99gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n665_), .B2(G99gat), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT112), .B(new_n664_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(G99gat), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT110), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n665_), .A2(new_n666_), .A3(G99gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n663_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n661_), .A2(KEYINPUT51), .ZN(new_n674_));
  AOI22_X1  g473(.A1(new_n661_), .A2(new_n669_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT51), .B1(new_n673_), .B2(KEYINPUT112), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n660_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT51), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n669_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT111), .B1(new_n673_), .B2(KEYINPUT112), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n664_), .B(new_n674_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT113), .B(new_n679_), .C1(new_n680_), .C2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n677_), .A2(new_n683_), .ZN(G1338gat));
  NAND3_X1  g483(.A1(new_n576_), .A2(new_n286_), .A3(new_n650_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G106gat), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT114), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT114), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n685_), .A2(new_n688_), .A3(G106gat), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT52), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n620_), .A2(new_n393_), .A3(new_n286_), .A4(new_n581_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n687_), .A2(KEYINPUT52), .A3(new_n689_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT53), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT53), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n692_), .A2(new_n697_), .A3(new_n693_), .A4(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1339gat));
  OAI211_X1 g498(.A(new_n491_), .B(new_n505_), .C1(new_n460_), .C2(new_n462_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT115), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n701_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n527_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT54), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n567_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT54), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT116), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n442_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT55), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT117), .ZN(new_n714_));
  INV_X1    g513(.A(new_n434_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n410_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n382_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n380_), .B1(new_n410_), .B2(new_n431_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(KEYINPUT12), .B2(new_n436_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n714_), .B(new_n444_), .C1(new_n717_), .C2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n444_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT117), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT55), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n442_), .A2(new_n711_), .A3(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n713_), .A2(new_n720_), .A3(new_n722_), .A4(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n450_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT56), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n728_), .A3(new_n450_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n727_), .A2(new_n490_), .A3(new_n456_), .A4(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n478_), .A2(new_n482_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n481_), .A2(new_n479_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n487_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT118), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n734_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n488_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n459_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n730_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n526_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT57), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT119), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n727_), .A2(new_n456_), .A3(new_n737_), .A4(new_n729_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT58), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n725_), .A2(new_n728_), .A3(new_n450_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n728_), .B1(new_n725_), .B2(new_n450_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n456_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n750_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n737_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n527_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n739_), .A2(KEYINPUT57), .A3(new_n526_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n742_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n566_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n710_), .A2(new_n756_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n370_), .A2(new_n583_), .A3(new_n236_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G113gat), .B1(new_n760_), .B2(new_n490_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT120), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT57), .B1(new_n739_), .B2(new_n526_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n526_), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n741_), .B(new_n764_), .C1(new_n730_), .C2(new_n738_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n762_), .B(new_n505_), .C1(new_n766_), .C2(new_n753_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT120), .B1(new_n755_), .B2(new_n566_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n710_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n758_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n770_), .A2(KEYINPUT59), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  AOI22_X1  g571(.A1(new_n706_), .A2(new_n709_), .B1(new_n755_), .B2(new_n566_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT59), .B1(new_n773_), .B2(new_n770_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n772_), .A2(new_n490_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n761_), .B1(new_n775_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g575(.A(KEYINPUT60), .ZN(new_n777_));
  XNOR2_X1  g576(.A(KEYINPUT121), .B(G120gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n532_), .B2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n757_), .A2(new_n758_), .A3(new_n779_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n772_), .A2(new_n463_), .A3(new_n774_), .A4(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n778_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n780_), .B2(KEYINPUT60), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT122), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n781_), .A2(KEYINPUT122), .A3(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(G1341gat));
  INV_X1    g587(.A(G127gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n759_), .B2(new_n566_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n790_), .A2(KEYINPUT123), .ZN(new_n791_));
  AND4_X1   g590(.A1(G127gat), .A2(new_n772_), .A3(new_n505_), .A4(new_n774_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n790_), .A2(KEYINPUT123), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(G1342gat));
  AOI21_X1  g593(.A(G134gat), .B1(new_n760_), .B2(new_n764_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n772_), .A2(G134gat), .A3(new_n774_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n567_), .ZN(G1343gat));
  AOI21_X1  g596(.A(new_n235_), .B1(new_n710_), .B2(new_n756_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n591_), .A2(new_n583_), .A3(new_n285_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n490_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n463_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(G148gat), .ZN(G1345gat));
  XOR2_X1   g604(.A(KEYINPUT124), .B(KEYINPUT125), .Z(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n800_), .B2(new_n566_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n806_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n798_), .A2(new_n505_), .A3(new_n799_), .A4(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT61), .B(G155gat), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n807_), .A2(new_n811_), .A3(new_n809_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1346gat));
  AOI21_X1  g614(.A(G162gat), .B1(new_n801_), .B2(new_n764_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n567_), .A2(G162gat), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT126), .Z(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n801_), .B2(new_n818_), .ZN(G1347gat));
  NOR2_X1   g618(.A1(new_n592_), .A2(new_n367_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n769_), .A2(new_n490_), .A3(new_n285_), .A4(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G169gat), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT62), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n769_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n286_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n826_), .A2(new_n490_), .A3(new_n223_), .A4(new_n820_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n821_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n824_), .A2(new_n827_), .A3(new_n828_), .ZN(G1348gat));
  NAND4_X1  g628(.A1(new_n769_), .A2(new_n463_), .A3(new_n285_), .A4(new_n820_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n208_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n773_), .A2(new_n286_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n832_), .A2(G176gat), .A3(new_n463_), .A4(new_n820_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT127), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT127), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n831_), .A2(new_n836_), .A3(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(G1349gat));
  INV_X1    g637(.A(new_n820_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n839_), .A2(new_n566_), .A3(new_n217_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n832_), .A2(new_n505_), .A3(new_n820_), .ZN(new_n841_));
  INV_X1    g640(.A(G183gat), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n826_), .A2(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(G1350gat));
  NAND4_X1  g642(.A1(new_n826_), .A2(new_n764_), .A3(new_n316_), .A4(new_n820_), .ZN(new_n844_));
  NOR4_X1   g643(.A1(new_n825_), .A2(new_n286_), .A3(new_n527_), .A4(new_n839_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n218_), .B2(new_n845_), .ZN(G1351gat));
  NOR2_X1   g645(.A1(new_n310_), .A2(new_n285_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n798_), .A2(new_n847_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n848_), .A2(new_n491_), .A3(new_n592_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(new_n256_), .ZN(G1352gat));
  NAND4_X1  g649(.A1(new_n798_), .A2(new_n463_), .A3(new_n847_), .A4(new_n591_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g651(.A1(new_n798_), .A2(new_n505_), .A3(new_n847_), .A4(new_n591_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n854_));
  AND2_X1   g653(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n853_), .B2(new_n854_), .ZN(G1354gat));
  INV_X1    g656(.A(G218gat), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n848_), .A2(new_n858_), .A3(new_n592_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n798_), .A2(new_n764_), .A3(new_n847_), .A4(new_n591_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n859_), .A2(new_n567_), .B1(new_n858_), .B2(new_n860_), .ZN(G1355gat));
endmodule


