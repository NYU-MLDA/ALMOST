//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n599_, new_n600_,
    new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n851_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G15gat), .B(G43gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT22), .B(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT74), .Z(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(G183gat), .B2(G190gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n211_), .A3(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n218_), .A2(new_n213_), .ZN(new_n219_));
  OR2_X1    g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n219_), .B(new_n221_), .C1(KEYINPUT24), .C2(new_n220_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n215_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT75), .B(KEYINPUT30), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n225_), .A2(KEYINPUT76), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(KEYINPUT76), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n206_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n206_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G127gat), .B(G134gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G113gat), .B(G120gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT77), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT31), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT78), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n229_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n234_), .A2(new_n235_), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n228_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n238_), .B1(new_n228_), .B2(new_n237_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G1gat), .B(G29gat), .ZN(new_n242_));
  INV_X1    g041(.A(G85gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT0), .B(G57gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  NAND2_X1  g045(.A1(G225gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT92), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G155gat), .A2(G162gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT79), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n252_), .B1(G155gat), .B2(G162gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(G141gat), .A2(G148gat), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(KEYINPUT3), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(KEYINPUT3), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G141gat), .A2(G148gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n255_), .A2(new_n256_), .A3(new_n259_), .A4(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n253_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT1), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n254_), .B(new_n257_), .C1(new_n252_), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(new_n233_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n232_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n249_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OR3_X1    g069(.A1(new_n267_), .A2(new_n233_), .A3(KEYINPUT93), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n267_), .A2(new_n233_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT93), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n249_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n248_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n268_), .A2(new_n269_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n247_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n246_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n246_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n270_), .A2(new_n271_), .B1(new_n249_), .B2(new_n274_), .ZN(new_n282_));
  OAI221_X1 g081(.A(new_n281_), .B1(new_n277_), .B2(new_n278_), .C1(new_n282_), .C2(new_n248_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n241_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286_));
  INV_X1    g085(.A(G92gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT18), .B(G64gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  XNOR2_X1  g089(.A(G197gat), .B(G204gat), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n291_), .A2(KEYINPUT86), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(KEYINPUT86), .ZN(new_n293_));
  XOR2_X1   g092(.A(G211gat), .B(G218gat), .Z(new_n294_));
  NAND4_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT21), .A4(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G204gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(KEYINPUT83), .A3(G197gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT21), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(new_n291_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT84), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT85), .B(KEYINPUT21), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n294_), .B1(new_n291_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n300_), .A2(new_n301_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n295_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(new_n220_), .A3(new_n211_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n219_), .B(new_n309_), .C1(new_n220_), .C2(new_n308_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n214_), .A2(new_n211_), .A3(new_n209_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT20), .B1(new_n307_), .B2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n307_), .A2(KEYINPUT87), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n307_), .A2(KEYINPUT87), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n313_), .B1(new_n316_), .B2(new_n223_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G226gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT91), .ZN(new_n322_));
  INV_X1    g121(.A(new_n223_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n314_), .A2(new_n323_), .A3(new_n315_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n320_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n321_), .B1(new_n322_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n322_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n290_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n327_), .A2(new_n322_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n290_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(new_n329_), .A4(new_n321_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT80), .B(KEYINPUT28), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT87), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n307_), .B(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n266_), .A2(KEYINPUT29), .ZN(new_n341_));
  NAND2_X1  g140(.A1(KEYINPUT81), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(KEYINPUT81), .A2(G233gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(G228gat), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT82), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n340_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT88), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n341_), .A2(new_n307_), .ZN(new_n350_));
  OAI22_X1  g149(.A1(new_n348_), .A2(new_n349_), .B1(new_n345_), .B2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n316_), .A2(new_n341_), .A3(new_n346_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(KEYINPUT88), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n338_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n350_), .A2(new_n345_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n352_), .B2(KEYINPUT88), .ZN(new_n356_));
  INV_X1    g155(.A(new_n338_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n348_), .A2(new_n349_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n266_), .A2(KEYINPUT29), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G78gat), .B(G106gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G22gat), .B(G50gat), .Z(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  AND3_X1   g163(.A1(new_n354_), .A2(new_n359_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n324_), .A2(new_n320_), .A3(new_n326_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n320_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n340_), .A2(new_n323_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n313_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n368_), .B1(new_n371_), .B2(KEYINPUT95), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n317_), .A2(new_n320_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT95), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n290_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(KEYINPUT27), .A3(new_n334_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n337_), .A2(new_n367_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT96), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n334_), .A2(KEYINPUT27), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n381_), .A2(new_n376_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT96), .B1(new_n382_), .B2(new_n367_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n285_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(KEYINPUT32), .B(new_n333_), .C1(new_n372_), .C2(new_n375_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n333_), .A2(KEYINPUT32), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n332_), .A2(new_n329_), .A3(new_n321_), .A4(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n284_), .A3(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n276_), .A2(new_n279_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT94), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(KEYINPUT33), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(new_n281_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n283_), .A2(new_n391_), .ZN(new_n394_));
  OAI221_X1 g193(.A(new_n246_), .B1(new_n277_), .B2(new_n248_), .C1(new_n282_), .C2(new_n278_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n388_), .B1(new_n396_), .B2(new_n335_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n367_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n365_), .A2(new_n366_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n284_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n337_), .A3(new_n377_), .A4(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n241_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n384_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT13), .ZN(new_n405_));
  XOR2_X1   g204(.A(KEYINPUT10), .B(G99gat), .Z(new_n406_));
  XOR2_X1   g205(.A(KEYINPUT64), .B(G106gat), .Z(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G85gat), .B(G92gat), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT9), .ZN(new_n410_));
  OR3_X1    g209(.A1(new_n243_), .A2(new_n287_), .A3(KEYINPUT9), .ZN(new_n411_));
  AND3_X1   g210(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .A4(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT8), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G99gat), .A2(G106gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n420_));
  NOR3_X1   g219(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT7), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n419_), .B(new_n420_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(KEYINPUT65), .A2(G99gat), .ZN(new_n424_));
  INV_X1    g223(.A(G106gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(KEYINPUT7), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n416_), .B(new_n409_), .C1(new_n423_), .C2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(KEYINPUT7), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n421_), .A2(new_n422_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n414_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n416_), .B1(new_n432_), .B2(new_n409_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n415_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT66), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT66), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n436_), .B(new_n415_), .C1(new_n429_), .C2(new_n433_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G57gat), .B(G64gat), .Z(new_n439_));
  INV_X1    g238(.A(KEYINPUT11), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G57gat), .B(G64gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n443_));
  XOR2_X1   g242(.A(G71gat), .B(G78gat), .Z(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n443_), .A2(new_n444_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n438_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  INV_X1    g248(.A(new_n447_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n435_), .A2(new_n450_), .A3(new_n437_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n438_), .A2(KEYINPUT67), .A3(new_n447_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n452_), .A2(G230gat), .A3(G233gat), .A4(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n447_), .A2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n434_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n438_), .B2(new_n447_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G230gat), .A2(G233gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n451_), .A2(new_n455_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G120gat), .B(G148gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(new_n296_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT5), .B(G176gat), .ZN(new_n464_));
  XOR2_X1   g263(.A(new_n463_), .B(new_n464_), .Z(new_n465_));
  NAND3_X1  g264(.A1(new_n454_), .A2(new_n461_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n454_), .B2(new_n461_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n405_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(KEYINPUT13), .A3(new_n466_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G29gat), .B(G36gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G43gat), .B(G50gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(G29gat), .B(G36gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT15), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT70), .B(G15gat), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(G22gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT70), .B(G15gat), .ZN(new_n484_));
  INV_X1    g283(.A(G22gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G1gat), .ZN(new_n487_));
  INV_X1    g286(.A(G8gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(new_n486_), .A3(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G1gat), .B(G8gat), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n483_), .A2(new_n491_), .A3(new_n486_), .A4(new_n489_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n481_), .A2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n475_), .A2(new_n478_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT71), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT71), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n479_), .A2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n498_), .A2(new_n493_), .A3(new_n494_), .A4(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT72), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT72), .B1(new_n481_), .B2(new_n495_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n498_), .A2(new_n500_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n495_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n501_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n504_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G113gat), .B(G141gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G169gat), .B(G197gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n507_), .B(new_n512_), .C1(KEYINPUT73), .C2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(KEYINPUT73), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT72), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(new_n496_), .B2(new_n501_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n520_), .A2(new_n511_), .A3(new_n505_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n512_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n518_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n472_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n404_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n438_), .A2(new_n497_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT34), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n530_), .A2(KEYINPUT35), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n481_), .B2(new_n434_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT69), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(KEYINPUT35), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT68), .Z(new_n535_));
  AOI22_X1  g334(.A1(new_n528_), .A2(new_n532_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n533_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n535_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n528_), .A2(KEYINPUT69), .A3(new_n540_), .A4(new_n532_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n545_), .B(KEYINPUT36), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n539_), .A2(new_n541_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT37), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n548_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n495_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(new_n447_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G127gat), .B(G155gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(G211gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT16), .B(G183gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT17), .Z(new_n563_));
  AND2_X1   g362(.A1(new_n558_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(KEYINPUT17), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n558_), .A2(new_n565_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n555_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n527_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n487_), .A3(new_n284_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT97), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT38), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n573_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n551_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(new_n567_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n527_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G1gat), .B1(new_n578_), .B2(new_n400_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(new_n575_), .A3(new_n579_), .ZN(G1324gat));
  OAI21_X1  g379(.A(G8gat), .B1(new_n578_), .B2(new_n382_), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT98), .B(KEYINPUT39), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n583_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n382_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n570_), .A2(new_n488_), .A3(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n584_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(G1325gat));
  OAI21_X1  g389(.A(G15gat), .B1(new_n578_), .B2(new_n241_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT100), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT41), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n569_), .A2(G15gat), .A3(new_n241_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT101), .Z(new_n597_));
  NAND3_X1  g396(.A1(new_n594_), .A2(new_n595_), .A3(new_n597_), .ZN(G1326gat));
  OAI21_X1  g397(.A(G22gat), .B1(new_n578_), .B2(new_n367_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT42), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n570_), .A2(new_n485_), .A3(new_n399_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1327gat));
  NAND4_X1  g401(.A1(new_n404_), .A2(KEYINPUT103), .A3(KEYINPUT43), .A4(new_n555_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n285_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n378_), .A2(new_n379_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n382_), .A2(KEYINPUT96), .A3(new_n367_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n604_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n241_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n398_), .B2(new_n401_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n555_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(KEYINPUT103), .A2(KEYINPUT43), .ZN(new_n611_));
  NAND2_X1  g410(.A1(KEYINPUT103), .A2(KEYINPUT43), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n526_), .A2(new_n567_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT102), .Z(new_n615_));
  NAND3_X1  g414(.A1(new_n603_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(KEYINPUT44), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n603_), .A2(new_n613_), .A3(new_n620_), .A4(new_n615_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n284_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G29gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n567_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n551_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n404_), .A2(new_n526_), .A3(new_n625_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n400_), .A2(G29gat), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(G1328gat));
  INV_X1    g427(.A(KEYINPUT106), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT46), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(KEYINPUT46), .ZN(new_n632_));
  INV_X1    g431(.A(G36gat), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n586_), .A2(new_n633_), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n626_), .A2(KEYINPUT45), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT45), .B1(new_n626_), .B2(new_n634_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n619_), .A2(new_n586_), .A3(new_n621_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT105), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n633_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n619_), .A2(KEYINPUT105), .A3(new_n586_), .A4(new_n621_), .ZN(new_n642_));
  AOI211_X1 g441(.A(new_n631_), .B(new_n638_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n640_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(G36gat), .A3(new_n642_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n630_), .B1(new_n645_), .B2(new_n637_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n643_), .A2(new_n646_), .ZN(G1329gat));
  NAND4_X1  g446(.A1(new_n619_), .A2(G43gat), .A3(new_n608_), .A4(new_n621_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT107), .B(G43gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n649_), .B1(new_n626_), .B2(new_n241_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g451(.A1(new_n619_), .A2(new_n399_), .A3(new_n621_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n626_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n367_), .A2(G50gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT108), .ZN(new_n656_));
  AOI22_X1  g455(.A1(new_n653_), .A2(G50gat), .B1(new_n654_), .B2(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT109), .Z(G1331gat));
  INV_X1    g457(.A(new_n472_), .ZN(new_n659_));
  AOI211_X1 g458(.A(new_n524_), .B(new_n659_), .C1(new_n384_), .C2(new_n403_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n577_), .ZN(new_n661_));
  INV_X1    g460(.A(G57gat), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n400_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n284_), .A3(new_n568_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n662_), .B2(new_n664_), .ZN(G1332gat));
  OAI21_X1  g464(.A(G64gat), .B1(new_n661_), .B2(new_n382_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT48), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n660_), .A2(new_n568_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n382_), .A2(G64gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n668_), .B2(new_n669_), .ZN(G1333gat));
  OAI21_X1  g469(.A(G71gat), .B1(new_n661_), .B2(new_n241_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT49), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n241_), .A2(G71gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n668_), .B2(new_n673_), .ZN(G1334gat));
  OAI21_X1  g473(.A(G78gat), .B1(new_n661_), .B2(new_n367_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT50), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n367_), .A2(G78gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n668_), .B2(new_n677_), .ZN(G1335gat));
  NAND2_X1  g477(.A1(new_n660_), .A2(new_n625_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G85gat), .B1(new_n680_), .B2(new_n284_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n603_), .A2(new_n613_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT110), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n603_), .A2(new_n613_), .A3(KEYINPUT110), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n659_), .A2(new_n524_), .A3(new_n624_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n684_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n400_), .A2(new_n243_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n681_), .B1(new_n687_), .B2(new_n688_), .ZN(G1336gat));
  NOR3_X1   g488(.A1(new_n679_), .A2(G92gat), .A3(new_n382_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n586_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(G92gat), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AOI211_X1 g493(.A(KEYINPUT111), .B(new_n690_), .C1(new_n691_), .C2(G92gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1337gat));
  NAND2_X1  g495(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n608_), .A2(new_n406_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n679_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n687_), .A2(new_n608_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(G99gat), .ZN(new_n701_));
  NOR2_X1   g500(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n702_), .B(new_n699_), .C1(new_n700_), .C2(G99gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1338gat));
  INV_X1    g505(.A(KEYINPUT52), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n603_), .A2(new_n613_), .A3(new_n399_), .A4(new_n686_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT113), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(G106gat), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n708_), .B2(G106gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n712_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(KEYINPUT52), .A3(new_n710_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n680_), .A2(new_n407_), .A3(new_n399_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n713_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT53), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT53), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n713_), .A2(new_n715_), .A3(new_n719_), .A4(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1339gat));
  AOI21_X1  g520(.A(new_n241_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n466_), .A2(new_n524_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n459_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT55), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n461_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n458_), .A2(new_n460_), .A3(KEYINPUT55), .A4(new_n459_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n465_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT56), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT56), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n734_), .B(new_n465_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n726_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n503_), .A2(new_n511_), .A3(new_n506_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n510_), .A2(new_n504_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n515_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n516_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n740_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n516_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n515_), .B1(new_n507_), .B2(new_n512_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT115), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n747_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n736_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n724_), .B1(new_n749_), .B2(new_n551_), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n576_), .B(new_n723_), .C1(new_n736_), .C2(new_n748_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n454_), .A2(new_n461_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n743_), .A2(new_n746_), .B1(new_n753_), .B2(new_n465_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n754_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT117), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT58), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT58), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n755_), .A2(KEYINPUT117), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n555_), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n624_), .B1(new_n752_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n567_), .A2(new_n524_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT114), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n469_), .A2(new_n763_), .A3(new_n471_), .A4(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n555_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n762_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT54), .B(new_n555_), .C1(new_n765_), .C2(new_n767_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n284_), .B(new_n722_), .C1(new_n761_), .C2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G113gat), .B1(new_n774_), .B2(new_n524_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT59), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n731_), .A2(new_n732_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n734_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n731_), .A2(KEYINPUT56), .A3(new_n732_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n725_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AOI22_X1  g581(.A1(new_n470_), .A2(new_n466_), .B1(new_n743_), .B2(new_n746_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n551_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n723_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n749_), .A2(new_n551_), .A3(new_n724_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n755_), .A2(KEYINPUT117), .A3(new_n758_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n758_), .B1(new_n755_), .B2(KEYINPUT117), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n769_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n567_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n555_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(new_n762_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n400_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n794_), .A2(KEYINPUT118), .A3(KEYINPUT59), .A4(new_n722_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n778_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n778_), .A2(new_n795_), .A3(KEYINPUT119), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n524_), .A2(G113gat), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT120), .Z(new_n802_));
  AOI21_X1  g601(.A(new_n775_), .B1(new_n800_), .B2(new_n802_), .ZN(G1340gat));
  INV_X1    g602(.A(G120gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n659_), .B2(KEYINPUT60), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n774_), .B(new_n805_), .C1(KEYINPUT60), .C2(new_n804_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT121), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n659_), .B1(new_n778_), .B2(new_n795_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n804_), .ZN(G1341gat));
  INV_X1    g608(.A(G127gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n774_), .A2(new_n810_), .A3(new_n624_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n567_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n810_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT122), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n811_), .C1(new_n812_), .C2(new_n810_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1342gat));
  AOI21_X1  g616(.A(G134gat), .B1(new_n774_), .B2(new_n576_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n555_), .A2(G134gat), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n800_), .B2(new_n819_), .ZN(G1343gat));
  NAND4_X1  g619(.A1(new_n794_), .A2(new_n399_), .A3(new_n382_), .A4(new_n241_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(new_n525_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT123), .B(G141gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1344gat));
  INV_X1    g623(.A(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n472_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g626(.A1(new_n821_), .A2(KEYINPUT124), .A3(new_n567_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT124), .B1(new_n821_), .B2(new_n567_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT61), .B(G155gat), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n830_), .B(new_n831_), .Z(G1346gat));
  INV_X1    g631(.A(G162gat), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n821_), .A2(new_n833_), .A3(new_n769_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n825_), .A2(new_n576_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n833_), .B2(new_n835_), .ZN(G1347gat));
  AOI21_X1  g635(.A(new_n382_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n604_), .A2(new_n399_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n837_), .A2(new_n524_), .A3(new_n207_), .A4(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT125), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n838_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n525_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n837_), .A2(KEYINPUT125), .A3(new_n524_), .A4(new_n838_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(G169gat), .A3(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(KEYINPUT62), .B2(new_n844_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT126), .B1(new_n844_), .B2(KEYINPUT62), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n839_), .B1(new_n846_), .B2(new_n847_), .ZN(G1348gat));
  NOR2_X1   g647(.A1(new_n841_), .A2(new_n659_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(new_n208_), .ZN(G1349gat));
  NOR2_X1   g649(.A1(new_n841_), .A2(new_n567_), .ZN(new_n851_));
  MUX2_X1   g650(.A(G183gat), .B(new_n216_), .S(new_n851_), .Z(G1350gat));
  OAI21_X1  g651(.A(G190gat), .B1(new_n841_), .B2(new_n769_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n576_), .A2(new_n217_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n841_), .B2(new_n854_), .ZN(G1351gat));
  NOR3_X1   g654(.A1(new_n608_), .A2(new_n367_), .A3(new_n284_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n837_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n524_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g659(.A1(new_n857_), .A2(new_n659_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n296_), .ZN(G1353gat));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n624_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n864_));
  AND2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n863_), .B2(new_n864_), .ZN(G1354gat));
  AOI21_X1  g666(.A(G218gat), .B1(new_n858_), .B2(new_n576_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n555_), .A2(G218gat), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n869_), .B(KEYINPUT127), .Z(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n858_), .B2(new_n870_), .ZN(G1355gat));
endmodule


