//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n207_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT9), .ZN(new_n213_));
  XOR2_X1   g012(.A(G85gat), .B(G92gat), .Z(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(KEYINPUT9), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n210_), .B(new_n215_), .C1(G106gat), .C2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220_));
  AND2_X1   g019(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n209_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n224_));
  NAND2_X1  g023(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n208_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n220_), .B1(new_n223_), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n209_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n208_), .A3(new_n225_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(KEYINPUT67), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT65), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n227_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n219_), .B1(new_n235_), .B2(new_n214_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n214_), .A2(new_n219_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n237_), .B1(new_n210_), .B2(new_n234_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n218_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G29gat), .B(G36gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G43gat), .B(G50gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT15), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G232gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT34), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT35), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n218_), .B(new_n242_), .C1(new_n236_), .C2(new_n238_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n244_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n247_), .A2(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n252_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n244_), .A2(new_n254_), .A3(new_n249_), .A4(new_n250_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n206_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n253_), .A2(KEYINPUT72), .A3(new_n255_), .A4(new_n205_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT37), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n256_), .A2(KEYINPUT36), .A3(new_n204_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G57gat), .B(G64gat), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n266_), .A2(KEYINPUT11), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(KEYINPUT11), .ZN(new_n268_));
  XOR2_X1   g067(.A(G71gat), .B(G78gat), .Z(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n268_), .A2(new_n269_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G15gat), .B(G22gat), .ZN(new_n273_));
  INV_X1    g072(.A(G1gat), .ZN(new_n274_));
  INV_X1    g073(.A(G8gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT14), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G1gat), .B(G8gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n272_), .B(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G231gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G127gat), .B(G155gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT16), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G183gat), .B(G211gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT17), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n282_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n287_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n282_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n265_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT73), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n296_));
  INV_X1    g095(.A(new_n272_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n239_), .A2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n272_), .B(new_n218_), .C1(new_n236_), .C2(new_n238_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(KEYINPUT12), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n239_), .A2(new_n301_), .A3(new_n297_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G230gat), .ZN(new_n304_));
  INV_X1    g103(.A(G233gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G176gat), .B(G204gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT69), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G120gat), .B(G148gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n308_), .A2(new_n310_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(KEYINPUT70), .ZN(new_n318_));
  INV_X1    g117(.A(new_n315_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n314_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n306_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n324_), .B1(new_n325_), .B2(new_n309_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n317_), .A2(new_n326_), .A3(KEYINPUT13), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT13), .B1(new_n317_), .B2(new_n326_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n296_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT13), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n323_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n325_), .A2(new_n309_), .A3(new_n320_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(KEYINPUT71), .A3(new_n327_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT98), .ZN(new_n338_));
  XOR2_X1   g137(.A(G8gat), .B(G36gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G204gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT85), .B1(new_n348_), .B2(G197gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n350_));
  INV_X1    g149(.A(G197gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(G204gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT21), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(G197gat), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n349_), .A2(new_n352_), .A3(new_n353_), .A4(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n348_), .A2(G197gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n351_), .A2(G204gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT21), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT86), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT86), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n355_), .A2(new_n358_), .A3(new_n362_), .A4(new_n359_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n359_), .A2(new_n353_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n349_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT87), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(KEYINPUT22), .B(G169gat), .Z(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT90), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n382_), .B2(G176gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n384_));
  INV_X1    g183(.A(G169gat), .ZN(new_n385_));
  INV_X1    g184(.A(G176gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT24), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n376_), .A2(new_n378_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n371_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n387_), .A2(KEYINPUT24), .A3(new_n388_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT25), .B(G183gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT26), .B(G190gat), .Z(new_n396_));
  OAI221_X1 g195(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n383_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n367_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT87), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n370_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n371_), .B(KEYINPUT77), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT78), .ZN(new_n405_));
  OR3_X1    g204(.A1(new_n404_), .A2(new_n393_), .A3(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n405_), .B1(new_n404_), .B2(new_n393_), .ZN(new_n407_));
  INV_X1    g206(.A(G190gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT26), .B1(new_n408_), .B2(KEYINPUT75), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n408_), .A2(KEYINPUT26), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n394_), .B(new_n409_), .C1(new_n410_), .C2(KEYINPUT75), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n406_), .A2(new_n391_), .A3(new_n407_), .A4(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n379_), .B(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n385_), .B2(KEYINPUT22), .ZN(new_n416_));
  AOI21_X1  g215(.A(G176gat), .B1(new_n385_), .B2(KEYINPUT22), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT22), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n373_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT80), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n373_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n412_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n403_), .B1(new_n426_), .B2(new_n369_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n347_), .B1(new_n402_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT96), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n383_), .A2(new_n397_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n369_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n399_), .A2(new_n412_), .A3(new_n425_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(KEYINPUT20), .A3(new_n432_), .ZN(new_n433_));
  OAI22_X1  g232(.A1(new_n428_), .A2(new_n429_), .B1(new_n346_), .B2(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n428_), .A2(new_n429_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n343_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n426_), .B2(new_n369_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n399_), .A2(new_n383_), .A3(new_n397_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n347_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n431_), .A2(KEYINPUT20), .A3(new_n346_), .A4(new_n432_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n343_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(KEYINPUT97), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT27), .ZN(new_n446_));
  INV_X1    g245(.A(new_n442_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n346_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n444_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT97), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n446_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n436_), .A2(new_n445_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n441_), .A2(new_n442_), .A3(new_n343_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT92), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n449_), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n443_), .A2(KEYINPUT92), .A3(new_n444_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n446_), .A3(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G127gat), .B(G134gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G113gat), .B(G120gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT3), .ZN(new_n463_));
  INV_X1    g262(.A(G141gat), .ZN(new_n464_));
  INV_X1    g263(.A(G148gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G141gat), .A2(G148gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT2), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n466_), .A2(new_n469_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(KEYINPUT1), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT1), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(G155gat), .A3(G162gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n479_), .A3(new_n473_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G141gat), .B(G148gat), .Z(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n462_), .A2(new_n483_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n472_), .A2(new_n475_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n461_), .A2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n484_), .A2(KEYINPUT4), .A3(new_n486_), .ZN(new_n491_));
  OR3_X1    g290(.A1(new_n461_), .A2(new_n485_), .A3(KEYINPUT4), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n489_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G1gat), .B(G29gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G85gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n490_), .A2(new_n494_), .A3(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n487_), .A2(new_n489_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n488_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n499_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT88), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT29), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n485_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G228gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT84), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n399_), .A2(new_n400_), .ZN(new_n512_));
  AOI211_X1 g311(.A(KEYINPUT87), .B(new_n367_), .C1(new_n361_), .C2(new_n363_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n510_), .B1(new_n399_), .B2(new_n508_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n506_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G78gat), .B(G106gat), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n483_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT28), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n485_), .B2(new_n507_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n518_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT28), .B1(new_n483_), .B2(KEYINPUT29), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n485_), .A2(new_n520_), .A3(new_n507_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n518_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G22gat), .B(G50gat), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n527_), .B(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n514_), .A2(new_n506_), .A3(new_n515_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n517_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n527_), .B(new_n528_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n531_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n533_), .B1(new_n534_), .B2(new_n516_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G15gat), .B(G43gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT82), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT30), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G227gat), .A2(G233gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(G71gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(G99gat), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n412_), .A2(new_n425_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n412_), .B2(new_n425_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n539_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n426_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n412_), .A2(new_n425_), .A3(new_n542_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n538_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT83), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT83), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n545_), .A2(new_n549_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n461_), .B(KEYINPUT31), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n551_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n556_));
  AND4_X1   g355(.A1(new_n552_), .A2(new_n545_), .A3(new_n549_), .A4(new_n554_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n532_), .B(new_n535_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n532_), .A2(new_n535_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n554_), .B1(new_n550_), .B2(KEYINPUT83), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n557_), .B1(new_n560_), .B2(new_n553_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n505_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n455_), .A2(new_n456_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n500_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(KEYINPUT94), .A3(KEYINPUT33), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT33), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n567_), .B1(new_n504_), .B2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n493_), .A2(new_n489_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n484_), .A2(new_n489_), .A3(new_n486_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n500_), .A2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT33), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n504_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n566_), .A2(new_n569_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n564_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n444_), .A2(KEYINPUT32), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n443_), .A2(new_n578_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n505_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n559_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(new_n561_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n458_), .A2(new_n563_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n242_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n279_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n243_), .A2(new_n279_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n279_), .B(new_n587_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n589_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n590_), .A2(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT74), .ZN(new_n596_));
  XOR2_X1   g395(.A(G169gat), .B(G197gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n594_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n338_), .B1(new_n586_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n581_), .A2(new_n505_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n434_), .A2(new_n435_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(new_n579_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n575_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n585_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n505_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n559_), .A2(new_n561_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n559_), .A2(new_n561_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n607_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n452_), .A2(new_n457_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n606_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(KEYINPUT98), .A3(new_n599_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n337_), .B1(new_n601_), .B2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n295_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n274_), .A3(new_n505_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n617_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n260_), .A2(new_n262_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n586_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n621_), .A2(new_n293_), .A3(new_n336_), .A4(new_n599_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n607_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n618_), .A2(new_n619_), .A3(new_n623_), .ZN(G1324gat));
  OAI21_X1  g423(.A(G8gat), .B1(new_n622_), .B2(new_n458_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT39), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n615_), .A2(new_n275_), .A3(new_n611_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n628_), .B(new_n630_), .ZN(G1325gat));
  INV_X1    g430(.A(new_n561_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G15gat), .B1(new_n622_), .B2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT41), .Z(new_n634_));
  INV_X1    g433(.A(G15gat), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n615_), .A2(new_n635_), .A3(new_n561_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(G1326gat));
  OAI21_X1  g436(.A(G22gat), .B1(new_n622_), .B2(new_n559_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n559_), .A2(G22gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT101), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n615_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(G1327gat));
  AOI211_X1 g442(.A(new_n293_), .B(new_n600_), .C1(new_n330_), .C2(new_n335_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n586_), .A2(KEYINPUT43), .A3(new_n265_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n620_), .A2(KEYINPUT37), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n646_), .B1(new_n612_), .B2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n644_), .B1(new_n645_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT43), .B1(new_n586_), .B2(new_n265_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n612_), .A2(new_n646_), .A3(new_n649_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(KEYINPUT44), .A3(new_n644_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n653_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(G29gat), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n607_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n620_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n293_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n614_), .A2(new_n505_), .A3(new_n662_), .ZN(new_n663_));
  AOI22_X1  g462(.A1(new_n658_), .A2(new_n660_), .B1(new_n659_), .B2(new_n663_), .ZN(G1328gat));
  NOR2_X1   g463(.A1(new_n458_), .A2(G36gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n614_), .A2(new_n662_), .A3(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n666_), .B(new_n667_), .Z(new_n668_));
  NAND3_X1  g467(.A1(new_n653_), .A2(new_n611_), .A3(new_n657_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(new_n670_), .A3(G36gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(G36gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n668_), .B(KEYINPUT46), .C1(new_n671_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1329gat));
  NAND3_X1  g476(.A1(new_n658_), .A2(G43gat), .A3(new_n561_), .ZN(new_n678_));
  INV_X1    g477(.A(G43gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n614_), .A2(new_n662_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(new_n632_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(G1330gat));
  NAND3_X1  g483(.A1(new_n658_), .A2(G50gat), .A3(new_n584_), .ZN(new_n685_));
  INV_X1    g484(.A(G50gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n680_), .B2(new_n559_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(G1331gat));
  NOR2_X1   g489(.A1(new_n292_), .A2(new_n599_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n621_), .A2(new_n337_), .A3(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT107), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n607_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n612_), .A2(new_n600_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT106), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(new_n337_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n295_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n607_), .A2(G57gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n695_), .B1(new_n699_), .B2(new_n700_), .ZN(G1332gat));
  OAI21_X1  g500(.A(G64gat), .B1(new_n694_), .B2(new_n458_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(KEYINPUT48), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(KEYINPUT48), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n458_), .A2(G64gat), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT108), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n703_), .A2(new_n704_), .B1(new_n699_), .B2(new_n706_), .ZN(G1333gat));
  NAND2_X1  g506(.A1(new_n693_), .A2(new_n561_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT49), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G71gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G71gat), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n632_), .A2(G71gat), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n710_), .A2(new_n711_), .B1(new_n699_), .B2(new_n712_), .ZN(G1334gat));
  OR3_X1    g512(.A1(new_n699_), .A2(G78gat), .A3(new_n559_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G78gat), .B1(new_n694_), .B2(new_n559_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(KEYINPUT50), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(KEYINPUT50), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n714_), .B1(new_n716_), .B2(new_n717_), .ZN(G1335gat));
  NOR3_X1   g517(.A1(new_n336_), .A2(new_n293_), .A3(new_n599_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n656_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n607_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n697_), .A2(new_n337_), .A3(new_n662_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n505_), .A2(new_n211_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(G1336gat));
  OAI21_X1  g523(.A(G92gat), .B1(new_n720_), .B2(new_n458_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n611_), .A2(new_n212_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n722_), .B2(new_n726_), .ZN(G1337gat));
  NOR2_X1   g526(.A1(new_n632_), .A2(new_n217_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n722_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G99gat), .B1(new_n720_), .B2(new_n632_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT109), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(KEYINPUT109), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n730_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n735_), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n737_), .B(new_n730_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1338gat));
  NOR2_X1   g538(.A1(new_n559_), .A2(G106gat), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n698_), .A2(KEYINPUT111), .A3(new_n662_), .A4(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742_));
  INV_X1    g541(.A(new_n740_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n722_), .B2(new_n743_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n741_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(G106gat), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n656_), .A2(new_n719_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(new_n584_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT112), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n748_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT53), .B1(new_n745_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n741_), .A2(new_n744_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n748_), .A2(new_n752_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .A4(new_n750_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(new_n758_), .ZN(G1339gat));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760_));
  INV_X1    g559(.A(G113gat), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT59), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n594_), .A2(new_n598_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n598_), .B1(new_n592_), .B2(new_n589_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n591_), .A2(new_n588_), .A3(new_n593_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n763_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(new_n333_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n303_), .A2(KEYINPUT55), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n306_), .A2(KEYINPUT114), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n325_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n323_), .B1(new_n775_), .B2(new_n771_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n776_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT58), .B(new_n769_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT115), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n769_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  INV_X1    g583(.A(new_n773_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n775_), .B1(new_n308_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n303_), .A2(KEYINPUT55), .A3(new_n771_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n324_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n776_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(KEYINPUT58), .A4(new_n769_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n780_), .A2(new_n783_), .A3(new_n649_), .A4(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n317_), .A2(new_n599_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n768_), .B1(new_n317_), .B2(new_n326_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n661_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(KEYINPUT57), .B(new_n661_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n334_), .A2(new_n327_), .A3(new_n691_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n334_), .A2(KEYINPUT113), .A3(new_n327_), .A4(new_n691_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n265_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT54), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(new_n810_), .A3(new_n265_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n802_), .A2(new_n292_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n611_), .A2(new_n607_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n562_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n762_), .B1(new_n812_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n795_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n797_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT57), .B1(new_n821_), .B2(new_n661_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n801_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n293_), .B1(new_n824_), .B2(new_n794_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n811_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n810_), .B1(new_n807_), .B2(new_n265_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT59), .B(new_n815_), .C1(new_n825_), .C2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n817_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n761_), .B1(new_n830_), .B2(new_n599_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n812_), .A2(new_n816_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n599_), .A2(new_n761_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n760_), .B1(new_n831_), .B2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n600_), .B1(new_n817_), .B2(new_n829_), .ZN(new_n837_));
  OAI221_X1 g636(.A(KEYINPUT116), .B1(new_n833_), .B2(new_n834_), .C1(new_n837_), .C2(new_n761_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1340gat));
  NOR2_X1   g638(.A1(new_n336_), .A2(KEYINPUT60), .ZN(new_n840_));
  MUX2_X1   g639(.A(new_n840_), .B(KEYINPUT60), .S(G120gat), .Z(new_n841_));
  NAND2_X1  g640(.A1(new_n832_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n336_), .B1(new_n817_), .B2(new_n829_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n843_), .A2(KEYINPUT117), .ZN(new_n844_));
  OAI21_X1  g643(.A(G120gat), .B1(new_n843_), .B2(KEYINPUT117), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n842_), .B1(new_n844_), .B2(new_n845_), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n832_), .A2(new_n847_), .A3(new_n293_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n292_), .B1(new_n817_), .B2(new_n829_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1342gat));
  AOI21_X1  g649(.A(G134gat), .B1(new_n832_), .B2(new_n620_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n851_), .A2(KEYINPUT118), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(KEYINPUT118), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n649_), .A2(G134gat), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n852_), .A2(new_n853_), .B1(new_n830_), .B2(new_n854_), .ZN(G1343gat));
  NOR2_X1   g654(.A1(new_n812_), .A2(new_n558_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n813_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n600_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n464_), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n336_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n465_), .ZN(G1345gat));
  NAND3_X1  g660(.A1(new_n856_), .A2(new_n293_), .A3(new_n813_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  INV_X1    g663(.A(G162gat), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n856_), .A2(new_n865_), .A3(new_n620_), .A4(new_n813_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n802_), .A2(new_n292_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n809_), .A2(new_n811_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n609_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n870_), .A2(new_n265_), .A3(new_n814_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n866_), .B1(new_n871_), .B2(new_n865_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT119), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n866_), .B(new_n874_), .C1(new_n871_), .C2(new_n865_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1347gat));
  NAND2_X1  g675(.A1(new_n611_), .A2(new_n607_), .ZN(new_n877_));
  NOR4_X1   g676(.A1(new_n812_), .A2(new_n584_), .A3(new_n632_), .A4(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n600_), .A2(new_n382_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT120), .Z(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n599_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(G169gat), .ZN(new_n884_));
  AOI211_X1 g683(.A(KEYINPUT62), .B(new_n385_), .C1(new_n878_), .C2(new_n599_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n881_), .B1(new_n884_), .B2(new_n885_), .ZN(G1348gat));
  NAND2_X1  g685(.A1(new_n878_), .A2(new_n337_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g687(.A1(new_n877_), .A2(new_n632_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n293_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n869_), .A2(new_n395_), .A3(new_n559_), .A4(new_n891_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n812_), .A2(new_n584_), .A3(new_n890_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n892_), .B(KEYINPUT121), .C1(new_n893_), .C2(G183gat), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n896_), .A3(new_n395_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n894_), .A2(new_n895_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n894_), .B2(new_n897_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1350gat));
  INV_X1    g699(.A(new_n396_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n878_), .A2(new_n620_), .A3(new_n901_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n878_), .A2(new_n649_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n408_), .ZN(G1351gat));
  INV_X1    g703(.A(new_n877_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n856_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(G197gat), .B1(new_n907_), .B2(new_n599_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n856_), .A2(G197gat), .A3(new_n599_), .A4(new_n905_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n910_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n908_), .A2(new_n911_), .A3(new_n912_), .ZN(G1352gat));
  NOR2_X1   g712(.A1(new_n906_), .A2(new_n336_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT124), .B(G204gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1353gat));
  AOI21_X1  g715(.A(new_n292_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n907_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT125), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT126), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n918_), .B(new_n921_), .ZN(G1354gat));
  XNOR2_X1  g721(.A(KEYINPUT127), .B(G218gat), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n906_), .A2(new_n265_), .A3(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n907_), .A2(new_n620_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n923_), .ZN(G1355gat));
endmodule


