//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  OR2_X1    g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  AND2_X1   g003(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n203_), .B(new_n207_), .C1(new_n204_), .C2(new_n205_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G85gat), .B(G92gat), .Z(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT8), .B1(new_n209_), .B2(KEYINPUT67), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n218_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .A4(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n217_), .A2(new_n216_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT10), .B(G99gat), .Z(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n221_), .A2(new_n222_), .A3(new_n203_), .A4(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n208_), .B(new_n209_), .C1(KEYINPUT67), .C2(KEYINPUT8), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n212_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n230_));
  XOR2_X1   g029(.A(G71gat), .B(G78gat), .Z(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n231_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n228_), .A2(KEYINPUT12), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n228_), .A2(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n212_), .A2(new_n226_), .A3(new_n227_), .A4(KEYINPUT68), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n235_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n236_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G230gat), .A2(G233gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(new_n235_), .A3(new_n239_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT12), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(new_n243_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT71), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT71), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n242_), .A2(new_n249_), .A3(new_n246_), .A4(new_n243_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n243_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n240_), .A2(new_n253_), .A3(new_n241_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n244_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n252_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT70), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n259_), .B(new_n252_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n251_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G120gat), .B(G148gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT5), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(G176gat), .ZN(new_n264_));
  INV_X1    g063(.A(G204gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n251_), .A2(new_n258_), .A3(new_n260_), .A4(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n267_), .A2(KEYINPUT13), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT13), .B1(new_n267_), .B2(new_n269_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT100), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G127gat), .B(G134gat), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(G113gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(G113gat), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n277_), .A2(G120gat), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(G120gat), .B1(new_n277_), .B2(new_n278_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT31), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT82), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n283_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  INV_X1    g091(.A(G169gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT22), .ZN(new_n295_));
  INV_X1    g094(.A(G176gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(G169gat), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n291_), .A2(new_n292_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT25), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n299_), .A2(KEYINPUT79), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(KEYINPUT79), .ZN(new_n301_));
  OAI21_X1  g100(.A(G183gat), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT80), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(KEYINPUT80), .B(G183gat), .C1(new_n300_), .C2(new_n301_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G190gat), .ZN(new_n306_));
  INV_X1    g105(.A(G183gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT25), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT78), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .A4(new_n309_), .ZN(new_n310_));
  OR3_X1    g109(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT81), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT81), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n318_), .A3(new_n315_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n312_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n298_), .B1(new_n310_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT30), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n286_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n286_), .A2(new_n322_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G71gat), .B(G99gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G15gat), .B(G43gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  NOR2_X1   g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n286_), .B(new_n322_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n328_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n275_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n325_), .A2(new_n328_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n331_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(KEYINPUT83), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n265_), .A2(G197gat), .ZN(new_n338_));
  INV_X1    g137(.A(G197gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G204gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n340_), .A3(KEYINPUT88), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT21), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n340_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n346_), .A2(new_n342_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(KEYINPUT21), .A3(new_n342_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT84), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n351_), .B1(G141gat), .B2(G148gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(KEYINPUT84), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n356_), .B(KEYINPUT1), .Z(new_n357_));
  NOR3_X1   g156(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AOI211_X1 g160(.A(new_n350_), .B(new_n355_), .C1(new_n357_), .C2(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n359_), .A2(new_n360_), .B1(G155gat), .B2(G162gat), .ZN(new_n363_));
  INV_X1    g162(.A(G141gat), .ZN(new_n364_));
  INV_X1    g163(.A(G148gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT86), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n364_), .B(new_n365_), .C1(new_n366_), .C2(KEYINPUT3), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n368_), .B(KEYINPUT86), .C1(G141gat), .C2(G148gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(G141gat), .A2(G148gat), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n371_), .A2(KEYINPUT2), .B1(new_n366_), .B2(KEYINPUT3), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n351_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n353_), .A2(KEYINPUT84), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT2), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n363_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT87), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT2), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n372_), .A3(new_n370_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(KEYINPUT87), .A3(new_n363_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n362_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n349_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G228gat), .ZN(new_n387_));
  INV_X1    g186(.A(G233gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  OAI221_X1 g189(.A(new_n349_), .B1(new_n387_), .B2(new_n388_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G78gat), .B(G106gat), .Z(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT89), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT28), .B(G22gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G50gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n355_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(G141gat), .B2(G148gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n360_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n356_), .B1(new_n400_), .B2(new_n358_), .ZN(new_n401_));
  OAI22_X1  g200(.A1(new_n353_), .A2(new_n380_), .B1(new_n368_), .B2(KEYINPUT86), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n369_), .B2(new_n367_), .ZN(new_n403_));
  AOI211_X1 g202(.A(new_n378_), .B(new_n401_), .C1(new_n403_), .C2(new_n381_), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT87), .B1(new_n382_), .B2(new_n363_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n399_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n397_), .B1(new_n406_), .B2(KEYINPUT29), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n384_), .A2(new_n385_), .A3(new_n396_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n394_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT90), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n390_), .A2(new_n391_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(new_n392_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT90), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n394_), .A2(new_n415_), .A3(new_n410_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n412_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n413_), .B(new_n392_), .Z(new_n418_));
  AOI21_X1  g217(.A(new_n415_), .B1(new_n394_), .B2(new_n410_), .ZN(new_n419_));
  AOI211_X1 g218(.A(KEYINPUT90), .B(new_n409_), .C1(new_n393_), .C2(KEYINPUT89), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n422_));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G64gat), .B(G92gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT19), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n291_), .A2(new_n292_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n297_), .A2(new_n294_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT25), .B(G183gat), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n306_), .A2(new_n433_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n311_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n431_), .A2(new_n432_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n430_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n438_), .A2(KEYINPUT96), .B1(new_n321_), .B2(new_n437_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n438_), .A2(KEYINPUT96), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n429_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n310_), .A2(new_n320_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n431_), .A2(new_n432_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n437_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n434_), .A2(new_n435_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n430_), .B1(new_n349_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n429_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n444_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n427_), .B1(new_n441_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT27), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n321_), .A2(new_n437_), .ZN(new_n452_));
  OAI211_X1 g251(.A(KEYINPUT20), .B(new_n448_), .C1(new_n349_), .C2(new_n446_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n448_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n426_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n450_), .A2(new_n451_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n426_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT92), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n454_), .A2(new_n455_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n427_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT92), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n462_), .B(new_n426_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n457_), .B1(new_n451_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G225gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n281_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n406_), .A2(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n281_), .B(new_n399_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(KEYINPUT4), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT4), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n406_), .A2(new_n471_), .A3(new_n467_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n466_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n466_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n474_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G1gat), .B(G29gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G85gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT0), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n479_), .B(G57gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n476_), .B(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n417_), .A2(new_n421_), .A3(new_n465_), .A4(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT98), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n480_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(KEYINPUT93), .A3(new_n486_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n459_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n470_), .A2(new_n466_), .A3(new_n472_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT94), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n468_), .A2(new_n469_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n480_), .B1(new_n496_), .B2(new_n474_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n470_), .A2(KEYINPUT94), .A3(new_n466_), .A4(new_n472_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT33), .B(new_n480_), .C1(new_n473_), .C2(new_n475_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n492_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT95), .B1(new_n491_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n481_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n427_), .A2(KEYINPUT32), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n504_), .B1(new_n441_), .B2(new_n449_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT97), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n460_), .A2(new_n504_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n503_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n492_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n502_), .A2(new_n508_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n417_), .A2(new_n421_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n337_), .B1(new_n484_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n465_), .B(KEYINPUT99), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n334_), .A2(new_n335_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n513_), .A3(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(new_n503_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G15gat), .B(G22gat), .Z(new_n521_));
  NAND2_X1  g320(.A1(G1gat), .A2(G8gat), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(KEYINPUT14), .B2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n523_), .B(KEYINPUT76), .Z(new_n524_));
  XOR2_X1   g323(.A(G1gat), .B(G8gat), .Z(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G29gat), .B(G36gat), .ZN(new_n527_));
  INV_X1    g326(.A(G43gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(G50gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n526_), .B(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(G229gat), .A3(G233gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n526_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n531_), .B(KEYINPUT15), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n537_), .B(KEYINPUT77), .Z(new_n538_));
  INV_X1    g337(.A(new_n531_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n536_), .B(new_n538_), .C1(new_n534_), .C2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G113gat), .B(G141gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(new_n293_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(new_n339_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n274_), .B1(new_n520_), .B2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(KEYINPUT100), .B(new_n547_), .C1(new_n515_), .C2(new_n519_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n273_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n539_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n535_), .A2(new_n228_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G134gat), .ZN(new_n561_));
  INV_X1    g360(.A(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT74), .Z(new_n566_));
  INV_X1    g365(.A(KEYINPUT73), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n558_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(new_n552_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n558_), .A2(new_n567_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n554_), .A2(new_n555_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n559_), .B(new_n566_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n558_), .B2(new_n557_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n563_), .B(new_n564_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n573_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT75), .B1(new_n575_), .B2(new_n576_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT37), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT37), .ZN(new_n580_));
  OAI221_X1 g379(.A(new_n573_), .B1(KEYINPUT75), .B2(new_n580_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n235_), .B(new_n584_), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n526_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G127gat), .B(G155gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT16), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(new_n307_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(G211gat), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n590_), .A2(new_n591_), .ZN(new_n593_));
  OR3_X1    g392(.A1(new_n586_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n586_), .A2(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n583_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n551_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(G1gat), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n503_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT38), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n577_), .B(KEYINPUT102), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT103), .Z(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n520_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n596_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n272_), .A2(new_n547_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n607_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G1gat), .B1(new_n611_), .B2(new_n481_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n602_), .A2(new_n603_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n604_), .A2(new_n612_), .A3(new_n613_), .ZN(G1324gat));
  INV_X1    g413(.A(G8gat), .ZN(new_n615_));
  INV_X1    g414(.A(new_n516_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n600_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G8gat), .B1(new_n611_), .B2(new_n516_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT39), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g420(.A(new_n337_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G15gat), .B1(new_n611_), .B2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT41), .Z(new_n624_));
  INV_X1    g423(.A(G15gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n600_), .A2(new_n625_), .A3(new_n337_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(G1326gat));
  INV_X1    g426(.A(G22gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n513_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n600_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G22gat), .B1(new_n611_), .B2(new_n513_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT42), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(G1327gat));
  AND2_X1   g432(.A1(new_n512_), .A2(new_n513_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n482_), .B(KEYINPUT98), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n622_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n519_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(KEYINPUT105), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n515_), .B2(new_n519_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n579_), .A2(KEYINPUT106), .A3(new_n581_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT106), .B1(new_n579_), .B2(new_n581_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n638_), .A2(new_n640_), .A3(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n582_), .A2(KEYINPUT43), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n520_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(new_n596_), .A3(new_n610_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n609_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(KEYINPUT44), .A3(new_n596_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n481_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n605_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n608_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n636_), .A2(new_n637_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT100), .B1(new_n660_), .B2(new_n547_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n550_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n272_), .B(new_n659_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT107), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n549_), .A2(new_n550_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n272_), .A4(new_n659_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(G29gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n503_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n657_), .A2(new_n670_), .ZN(G1328gat));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  INV_X1    g471(.A(G36gat), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n664_), .A2(new_n673_), .A3(new_n616_), .A4(new_n667_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT45), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n653_), .A2(new_n616_), .A3(new_n655_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G36gat), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT108), .B(new_n672_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n668_), .A2(KEYINPUT45), .A3(new_n673_), .A4(new_n616_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n674_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT44), .B1(new_n654_), .B2(new_n596_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n648_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n683_));
  NOR4_X1   g482(.A1(new_n683_), .A2(new_n652_), .A3(new_n608_), .A4(new_n609_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n682_), .A2(new_n684_), .A3(new_n516_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n679_), .B(new_n681_), .C1(new_n685_), .C2(new_n673_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT46), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n678_), .A2(new_n688_), .ZN(G1329gat));
  INV_X1    g488(.A(new_n517_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G43gat), .B1(new_n656_), .B2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n668_), .A2(new_n528_), .A3(new_n337_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1330gat));
  OAI21_X1  g494(.A(G50gat), .B1(new_n656_), .B2(new_n513_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n668_), .A2(new_n530_), .A3(new_n629_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1331gat));
  NOR2_X1   g497(.A1(new_n272_), .A2(new_n547_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n607_), .A2(new_n608_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(G57gat), .A3(new_n503_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT110), .Z(new_n703_));
  NOR3_X1   g502(.A1(new_n520_), .A2(new_n547_), .A3(new_n272_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n597_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT109), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n481_), .B1(new_n705_), .B2(KEYINPUT109), .ZN(new_n707_));
  AOI21_X1  g506(.A(G57gat), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n703_), .A2(new_n708_), .ZN(G1332gat));
  OR3_X1    g508(.A1(new_n705_), .A2(G64gat), .A3(new_n516_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G64gat), .B1(new_n700_), .B2(new_n516_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT111), .Z(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(KEYINPUT48), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(KEYINPUT48), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(G1333gat));
  OR3_X1    g514(.A1(new_n705_), .A2(G71gat), .A3(new_n622_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G71gat), .B1(new_n700_), .B2(new_n622_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT112), .Z(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(KEYINPUT49), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(KEYINPUT49), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1334gat));
  OAI21_X1  g520(.A(G78gat), .B1(new_n700_), .B2(new_n513_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT50), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n513_), .A2(G78gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n705_), .B2(new_n724_), .ZN(G1335gat));
  NAND2_X1  g524(.A1(new_n704_), .A2(new_n659_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G85gat), .B1(new_n727_), .B2(new_n503_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n699_), .A2(new_n596_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n683_), .A2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n481_), .A2(new_n213_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n728_), .B1(new_n730_), .B2(new_n731_), .ZN(G1336gat));
  AOI21_X1  g531(.A(G92gat), .B1(new_n727_), .B2(new_n616_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n516_), .A2(new_n218_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n730_), .B2(new_n734_), .ZN(G1337gat));
  AND3_X1   g534(.A1(new_n727_), .A2(new_n517_), .A3(new_n223_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n730_), .A2(new_n337_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G99gat), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g538(.A1(new_n727_), .A2(new_n224_), .A3(new_n629_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n730_), .A2(new_n629_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(G106gat), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n683_), .A2(new_n513_), .A3(new_n729_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT113), .B1(new_n744_), .B2(new_n224_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n743_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n740_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n740_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1339gat));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n251_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n242_), .A2(new_n246_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n252_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n242_), .A2(KEYINPUT55), .A3(new_n246_), .A4(new_n243_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n755_), .A2(KEYINPUT116), .A3(new_n757_), .A4(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT55), .B1(new_n248_), .B2(new_n250_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n757_), .A2(new_n758_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n759_), .A2(new_n763_), .A3(new_n266_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT56), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n759_), .A2(new_n763_), .A3(new_n766_), .A4(new_n266_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n765_), .A2(new_n547_), .A3(new_n269_), .A4(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n267_), .A2(new_n269_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n532_), .A2(new_n538_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n536_), .B1(new_n534_), .B2(new_n539_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n770_), .B(new_n544_), .C1(new_n771_), .C2(new_n538_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n545_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n769_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n768_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n658_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n765_), .A2(new_n269_), .A3(new_n773_), .A4(new_n767_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n781_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n583_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n605_), .B1(new_n768_), .B2(new_n774_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT117), .B1(new_n785_), .B2(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(KEYINPUT57), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n779_), .A2(new_n784_), .A3(new_n786_), .A4(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n596_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n271_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n267_), .A2(KEYINPUT13), .A3(new_n269_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n790_), .A2(new_n608_), .A3(new_n548_), .A4(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n272_), .A2(KEYINPUT114), .A3(new_n608_), .A4(new_n548_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n582_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT115), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n794_), .A2(new_n795_), .A3(new_n798_), .A4(new_n582_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n797_), .A2(KEYINPUT54), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n799_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n789_), .A2(new_n800_), .A3(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n518_), .A2(new_n481_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G113gat), .B1(new_n807_), .B2(new_n547_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n776_), .A2(new_n778_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n784_), .A2(new_n809_), .A3(new_n787_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n803_), .B(new_n800_), .C1(new_n810_), .C2(new_n608_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n518_), .A2(KEYINPUT59), .A3(new_n481_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n806_), .A2(KEYINPUT59), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n547_), .A2(G113gat), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n808_), .B1(new_n813_), .B2(new_n814_), .ZN(G1340gat));
  INV_X1    g614(.A(G120gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n272_), .B2(KEYINPUT60), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT118), .B1(new_n816_), .B2(KEYINPUT60), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n806_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n813_), .A2(new_n273_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n821_), .B1(new_n823_), .B2(new_n816_), .ZN(G1341gat));
  NAND2_X1  g623(.A1(new_n803_), .A2(new_n800_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n596_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G127gat), .B1(new_n827_), .B2(new_n805_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n608_), .A2(G127gat), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT119), .Z(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n813_), .B2(new_n830_), .ZN(G1342gat));
  AOI21_X1  g630(.A(G134gat), .B1(new_n807_), .B2(new_n606_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n583_), .A2(G134gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n813_), .B2(new_n833_), .ZN(G1343gat));
  NOR4_X1   g633(.A1(new_n337_), .A2(new_n616_), .A3(new_n481_), .A4(new_n513_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n788_), .A2(new_n596_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n825_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT120), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n804_), .A2(new_n839_), .A3(new_n835_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n547_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n273_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n608_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  AND2_X1   g647(.A1(new_n606_), .A2(new_n562_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n804_), .A2(new_n839_), .A3(new_n835_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n839_), .B1(new_n804_), .B2(new_n835_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n643_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n854_), .B2(new_n562_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT121), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n852_), .B(new_n857_), .C1(new_n854_), .C2(new_n562_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1347gat));
  XOR2_X1   g658(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n860_));
  NOR4_X1   g659(.A1(new_n622_), .A2(new_n503_), .A3(new_n629_), .A4(new_n516_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n811_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n547_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n860_), .B1(new_n864_), .B2(KEYINPUT22), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n293_), .ZN(new_n866_));
  OAI211_X1 g665(.A(G169gat), .B(new_n860_), .C1(new_n864_), .C2(KEYINPUT22), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n866_), .B(new_n867_), .C1(new_n860_), .C2(new_n864_), .ZN(G1348gat));
  AND4_X1   g667(.A1(G176gat), .A2(new_n804_), .A3(new_n273_), .A4(new_n861_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n296_), .B1(new_n862_), .B2(new_n272_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n870_), .A2(KEYINPUT123), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(KEYINPUT123), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n871_), .B2(new_n872_), .ZN(G1349gat));
  AOI21_X1  g672(.A(G183gat), .B1(new_n827_), .B2(new_n861_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n862_), .A2(new_n596_), .A3(new_n433_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1350gat));
  OAI21_X1  g675(.A(G190gat), .B1(new_n862_), .B2(new_n582_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n606_), .A2(new_n306_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n862_), .B2(new_n878_), .ZN(G1351gat));
  AOI21_X1  g678(.A(new_n337_), .B1(new_n826_), .B2(new_n789_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n516_), .A2(new_n503_), .A3(new_n513_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n547_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n882_), .A2(new_n883_), .A3(new_n339_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n882_), .B2(new_n339_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n882_), .A2(new_n339_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(G1352gat));
  NAND2_X1  g686(.A1(new_n880_), .A2(new_n881_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n272_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n265_), .ZN(G1353gat));
  NAND2_X1  g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n880_), .A2(new_n608_), .A3(new_n881_), .A4(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  OR3_X1    g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n888_), .B2(new_n596_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n893_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(G1354gat));
  NAND4_X1  g697(.A1(new_n804_), .A2(new_n622_), .A3(new_n606_), .A4(new_n881_), .ZN(new_n899_));
  INV_X1    g698(.A(G218gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n583_), .A2(G218gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT126), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n888_), .B2(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


