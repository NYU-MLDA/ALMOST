//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n976_, new_n977_, new_n978_, new_n980_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n991_, new_n992_, new_n993_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  AOI22_X1  g011(.A1(new_n208_), .A2(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT26), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT26), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(G190gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n215_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n206_), .B(new_n213_), .C1(new_n218_), .C2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT77), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT22), .B1(new_n224_), .B2(new_n202_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT22), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G169gat), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n225_), .B(new_n203_), .C1(new_n224_), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n207_), .A2(new_n209_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n229_), .B(new_n230_), .C1(G183gat), .C2(G190gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n231_), .A3(new_n205_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n223_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT30), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(KEYINPUT79), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(KEYINPUT79), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT78), .B(G15gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G227gat), .A2(G233gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n235_), .A2(new_n236_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n236_), .A2(new_n243_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G127gat), .B(G134gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT31), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n245_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(new_n254_), .B2(new_n251_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(G85gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G57gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT81), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT81), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n268_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT3), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G141gat), .A2(G148gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n267_), .A2(new_n269_), .A3(new_n272_), .A4(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT82), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT82), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n279_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n265_), .B1(new_n276_), .B2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n283_), .A2(new_n273_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT1), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n263_), .A2(new_n286_), .A3(new_n264_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n282_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT83), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT83), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n282_), .A2(new_n291_), .A3(new_n288_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n292_), .A3(new_n250_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n289_), .A2(new_n250_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT4), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT4), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n290_), .A2(new_n298_), .A3(new_n292_), .A4(new_n250_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n295_), .A2(KEYINPUT96), .A3(new_n297_), .A4(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n293_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n297_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT96), .B1(new_n304_), .B2(new_n295_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n262_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT96), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n293_), .A2(KEYINPUT4), .A3(new_n294_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n307_), .B1(new_n308_), .B2(new_n303_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n309_), .A2(new_n261_), .A3(new_n301_), .A4(new_n300_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n306_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G8gat), .B(G36gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT32), .ZN(new_n317_));
  INV_X1    g116(.A(G197gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(G204gat), .ZN(new_n319_));
  INV_X1    g118(.A(G204gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT87), .B1(new_n320_), .B2(G197gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(new_n318_), .A3(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n319_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT21), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G211gat), .B(G218gat), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT86), .B1(new_n318_), .B2(G204gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT86), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(new_n320_), .A3(G197gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n318_), .A2(G204gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n328_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT21), .ZN(new_n333_));
  INV_X1    g132(.A(new_n326_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n334_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n327_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n202_), .A2(KEYINPUT22), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n227_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n231_), .B(new_n205_), .C1(G176gat), .C2(new_n338_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT91), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT91), .B1(new_n220_), .B2(new_n221_), .ZN(new_n341_));
  INV_X1    g140(.A(G183gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT25), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G183gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n340_), .A2(new_n341_), .A3(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n348_));
  NOR2_X1   g147(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n204_), .B(new_n205_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n349_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n212_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n208_), .A2(new_n210_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n347_), .A2(KEYINPUT93), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT93), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n350_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n220_), .A2(new_n221_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT91), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT91), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n214_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n357_), .B1(new_n358_), .B2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n336_), .B(new_n339_), .C1(new_n356_), .C2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT19), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  INV_X1    g168(.A(new_n319_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n322_), .B1(new_n318_), .B2(G204gat), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n320_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n325_), .B(new_n370_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n333_), .A2(new_n373_), .A3(new_n326_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(KEYINPUT21), .A3(new_n334_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n223_), .A2(new_n232_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n369_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n365_), .A2(new_n368_), .A3(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n374_), .A2(new_n376_), .A3(new_n223_), .A4(new_n232_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT20), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n339_), .B1(new_n356_), .B2(new_n364_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n383_), .B2(new_n377_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n380_), .B1(new_n384_), .B2(new_n368_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT97), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n317_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n339_), .B1(new_n347_), .B2(new_n355_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT98), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT98), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n390_), .B(new_n339_), .C1(new_n347_), .C2(new_n355_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n336_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n368_), .B1(new_n392_), .B2(new_n379_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT99), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n394_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n369_), .B1(new_n336_), .B2(new_n233_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n339_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT93), .B1(new_n347_), .B2(new_n355_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n358_), .A2(new_n357_), .A3(new_n363_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n397_), .B(new_n368_), .C1(new_n401_), .C2(new_n336_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n395_), .A2(new_n396_), .A3(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(KEYINPUT32), .B(new_n316_), .C1(new_n385_), .C2(KEYINPUT97), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n387_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n311_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT100), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT100), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n311_), .A2(new_n405_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n302_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n410_), .A2(KEYINPUT33), .A3(new_n261_), .A4(new_n309_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n316_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n385_), .A2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n397_), .B1(new_n401_), .B2(new_n336_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n367_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n380_), .A3(new_n316_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(KEYINPUT95), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT95), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n415_), .A2(new_n418_), .A3(new_n380_), .A4(new_n316_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n310_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n295_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n293_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n262_), .A3(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n411_), .A2(new_n420_), .A3(new_n422_), .A4(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n407_), .A2(new_n409_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G228gat), .ZN(new_n428_));
  OR2_X1    g227(.A1(KEYINPUT85), .A2(G233gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(KEYINPUT85), .A2(G233gat), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(new_n282_), .B2(new_n288_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n433_), .B2(new_n336_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n290_), .A2(KEYINPUT29), .A3(new_n292_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n336_), .A2(new_n431_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n435_), .A2(KEYINPUT88), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT88), .B1(new_n435_), .B2(new_n436_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n434_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G78gat), .B(G106gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n434_), .B(new_n440_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(G22gat), .B(G50gat), .Z(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n290_), .A2(new_n292_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n448_), .B1(new_n449_), .B2(new_n432_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n278_), .A2(new_n280_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n270_), .A2(new_n271_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n451_), .A2(new_n269_), .A3(new_n452_), .A4(new_n267_), .ZN(new_n453_));
  AOI221_X4 g252(.A(KEYINPUT83), .B1(new_n287_), .B2(new_n285_), .C1(new_n453_), .C2(new_n265_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n291_), .B1(new_n282_), .B2(new_n288_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n432_), .B(new_n448_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n446_), .B1(new_n450_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n432_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n447_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n445_), .A3(new_n456_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT90), .B1(new_n444_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n466_));
  AOI211_X1 g265(.A(new_n466_), .B(new_n462_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n442_), .A2(new_n462_), .A3(new_n443_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n442_), .A2(KEYINPUT89), .A3(new_n462_), .A4(new_n443_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n465_), .A2(new_n468_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n427_), .A2(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n469_), .A2(new_n470_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n472_), .ZN(new_n476_));
  OAI22_X1  g275(.A1(new_n475_), .A2(new_n476_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT27), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n417_), .A2(new_n478_), .A3(new_n419_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT103), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n417_), .A2(KEYINPUT103), .A3(new_n478_), .A4(new_n419_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n402_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n483_));
  AOI211_X1 g282(.A(KEYINPUT99), .B(new_n368_), .C1(new_n392_), .C2(new_n379_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n412_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT101), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(KEYINPUT101), .B(new_n412_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n478_), .B1(new_n416_), .B2(KEYINPUT102), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT102), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n415_), .A2(new_n491_), .A3(new_n380_), .A4(new_n316_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n481_), .A2(new_n482_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n311_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n477_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n257_), .B1(new_n474_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n494_), .ZN(new_n498_));
  NOR4_X1   g297(.A1(new_n498_), .A2(new_n477_), .A3(new_n256_), .A4(new_n311_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G169gat), .B(G197gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G15gat), .B(G22gat), .ZN(new_n505_));
  INV_X1    g304(.A(G1gat), .ZN(new_n506_));
  INV_X1    g305(.A(G8gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G1gat), .B(G8gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  XNOR2_X1  g310(.A(G29gat), .B(G36gat), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n512_), .A2(KEYINPUT71), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(KEYINPUT71), .ZN(new_n514_));
  XOR2_X1   g313(.A(G43gat), .B(G50gat), .Z(new_n515_));
  OR3_X1    g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n515_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n511_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n517_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT15), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n516_), .A2(new_n517_), .A3(KEYINPUT15), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n509_), .B(new_n510_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n520_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n521_), .A2(new_n526_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n519_), .B1(new_n528_), .B2(new_n518_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n504_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n524_), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT15), .B1(new_n516_), .B2(new_n517_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n526_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n520_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n529_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT75), .B1(new_n535_), .B2(new_n503_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT75), .ZN(new_n537_));
  NOR4_X1   g336(.A1(new_n527_), .A2(new_n537_), .A3(new_n529_), .A4(new_n504_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n530_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n500_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(G85gat), .ZN(new_n544_));
  INV_X1    g343(.A(G92gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT6), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT6), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(G99gat), .A3(G106gat), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT7), .ZN(new_n555_));
  INV_X1    g354(.A(G99gat), .ZN(new_n556_));
  INV_X1    g355(.A(G106gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n549_), .B1(new_n554_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT8), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(KEYINPUT67), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n551_), .A2(new_n553_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(new_n559_), .A3(new_n558_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(new_n549_), .A3(new_n563_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT10), .B(G99gat), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT65), .B1(new_n570_), .B2(G106gat), .ZN(new_n571_));
  OR2_X1    g370(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT65), .ZN(new_n573_));
  NAND2_X1  g372(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n557_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n546_), .A2(KEYINPUT9), .A3(new_n547_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n547_), .A2(KEYINPUT9), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n577_), .A2(new_n566_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT66), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT66), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n576_), .A2(new_n582_), .A3(new_n579_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n569_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT11), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT11), .ZN(new_n587_));
  XOR2_X1   g386(.A(G71gat), .B(G78gat), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n543_), .B1(new_n584_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT64), .Z(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n559_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AOI211_X1 g397(.A(new_n548_), .B(new_n564_), .C1(new_n598_), .C2(new_n566_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n563_), .B1(new_n567_), .B2(new_n549_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n576_), .A2(new_n582_), .A3(new_n579_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n582_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n601_), .B(new_n591_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n601_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n591_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(KEYINPUT12), .A3(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n592_), .A2(new_n595_), .A3(new_n604_), .A4(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT69), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n542_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n604_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT69), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n595_), .A4(new_n607_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n581_), .A2(new_n583_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n591_), .B1(new_n615_), .B2(new_n601_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n594_), .B1(new_n616_), .B2(new_n611_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n609_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT5), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n620_), .B(new_n621_), .Z(new_n622_));
  NAND2_X1  g421(.A1(new_n618_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n609_), .A2(new_n614_), .A3(new_n617_), .A4(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n626_), .A2(KEYINPUT13), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(KEYINPUT13), .A3(new_n625_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT70), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT70), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n584_), .A2(new_n521_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n636_), .B1(new_n525_), .B2(new_n584_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT34), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(KEYINPUT35), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n640_), .A2(KEYINPUT35), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n642_), .A2(KEYINPUT72), .B1(new_n637_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT72), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n638_), .A2(new_n646_), .A3(new_n641_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(G134gat), .B(G162gat), .Z(new_n649_));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT36), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n648_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n645_), .A2(new_n652_), .A3(new_n651_), .A4(new_n647_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT37), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n655_), .A2(KEYINPUT37), .A3(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(G231gat), .A2(G233gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n526_), .B(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(new_n606_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT74), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  XOR2_X1   g465(.A(G127gat), .B(G155gat), .Z(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(G183gat), .B(G211gat), .Z(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT17), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n666_), .B(new_n672_), .ZN(new_n673_));
  OR3_X1    g472(.A1(new_n664_), .A2(KEYINPUT17), .A3(new_n671_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n661_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n541_), .A2(new_n635_), .A3(new_n677_), .ZN(new_n678_));
  OR3_X1    g477(.A1(new_n678_), .A2(G1gat), .A3(new_n495_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT38), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n657_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n500_), .A2(new_n682_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n683_), .A2(new_n539_), .A3(new_n635_), .A4(new_n675_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G1gat), .B1(new_n684_), .B2(new_n495_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(new_n680_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n681_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT104), .ZN(G1324gat));
  NOR3_X1   g487(.A1(new_n678_), .A2(G8gat), .A3(new_n494_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G8gat), .B1(new_n684_), .B2(new_n494_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n690_), .A2(KEYINPUT39), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(KEYINPUT39), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n693_), .B(new_n695_), .ZN(G1325gat));
  OAI21_X1  g495(.A(G15gat), .B1(new_n684_), .B2(new_n256_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT41), .Z(new_n698_));
  OR2_X1    g497(.A1(new_n256_), .A2(G15gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n678_), .B2(new_n699_), .ZN(G1326gat));
  OAI21_X1  g499(.A(G22gat), .B1(new_n684_), .B2(new_n473_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT42), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n473_), .A2(G22gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n678_), .B2(new_n703_), .ZN(G1327gat));
  INV_X1    g503(.A(new_n661_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n420_), .A2(new_n422_), .A3(new_n425_), .ZN(new_n706_));
  AOI22_X1  g505(.A1(new_n706_), .A2(new_n411_), .B1(new_n406_), .B2(KEYINPUT100), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n477_), .B1(new_n707_), .B2(new_n409_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n477_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n256_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n498_), .A2(new_n477_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n256_), .A2(new_n311_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n705_), .B1(new_n710_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT107), .B(KEYINPUT43), .C1(new_n714_), .C2(new_n715_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n634_), .A2(new_n540_), .A3(new_n675_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n714_), .B2(KEYINPUT107), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n661_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(KEYINPUT106), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n716_), .B(new_n717_), .C1(new_n719_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT107), .B1(new_n714_), .B2(new_n715_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT43), .B1(new_n721_), .B2(new_n720_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n728_), .A2(KEYINPUT44), .A3(new_n716_), .A4(new_n717_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n725_), .A2(G29gat), .A3(new_n729_), .A4(new_n311_), .ZN(new_n730_));
  INV_X1    g529(.A(G29gat), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n657_), .A2(new_n675_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n541_), .A2(new_n635_), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n733_), .B2(new_n495_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n725_), .A2(new_n498_), .A3(new_n729_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G36gat), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n494_), .A2(G36gat), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n733_), .A2(new_n738_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT45), .Z(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n737_), .A2(KEYINPUT46), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1329gat));
  NAND4_X1  g544(.A1(new_n725_), .A2(G43gat), .A3(new_n257_), .A4(new_n729_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n238_), .B1(new_n733_), .B2(new_n256_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g548(.A1(new_n733_), .A2(G50gat), .A3(new_n473_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n725_), .A2(new_n477_), .A3(new_n729_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(KEYINPUT108), .ZN(new_n752_));
  OAI21_X1  g551(.A(G50gat), .B1(new_n751_), .B2(KEYINPUT108), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(G1331gat));
  NAND2_X1  g553(.A1(new_n675_), .A2(new_n540_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n635_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n683_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G57gat), .B1(new_n757_), .B2(new_n495_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n634_), .A2(new_n677_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT109), .Z(new_n760_));
  NOR2_X1   g559(.A1(new_n500_), .A2(new_n539_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n495_), .A2(G57gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n758_), .B1(new_n763_), .B2(new_n764_), .ZN(G1332gat));
  INV_X1    g564(.A(G64gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n766_), .A3(new_n498_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n757_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n768_), .B2(new_n498_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT48), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n769_), .A2(new_n770_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n767_), .B1(new_n772_), .B2(new_n773_), .ZN(G1333gat));
  OAI21_X1  g573(.A(G71gat), .B1(new_n757_), .B2(new_n256_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT49), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n256_), .A2(G71gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n763_), .B2(new_n777_), .ZN(G1334gat));
  OAI21_X1  g577(.A(G78gat), .B1(new_n757_), .B2(new_n473_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT50), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n473_), .A2(G78gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n763_), .B2(new_n781_), .ZN(G1335gat));
  AND2_X1   g581(.A1(new_n728_), .A2(new_n716_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n635_), .A2(new_n539_), .A3(new_n675_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n544_), .B1(new_n785_), .B2(new_n311_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n634_), .A2(new_n732_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n761_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n788_), .A2(G85gat), .A3(new_n495_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n786_), .A2(new_n789_), .ZN(G1336gat));
  AOI21_X1  g589(.A(new_n545_), .B1(new_n785_), .B2(new_n498_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n788_), .A2(G92gat), .A3(new_n494_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1337gat));
  NAND3_X1  g592(.A1(new_n783_), .A2(new_n257_), .A3(new_n784_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G99gat), .ZN(new_n795_));
  OR3_X1    g594(.A1(new_n788_), .A2(new_n256_), .A3(new_n570_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT51), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(new_n799_), .A3(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1338gat));
  NAND4_X1  g600(.A1(new_n787_), .A2(new_n761_), .A3(new_n557_), .A4(new_n477_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n728_), .A2(new_n477_), .A3(new_n716_), .A4(new_n784_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n803_), .A2(new_n804_), .A3(G106gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n803_), .B2(G106gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT53), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n802_), .B(new_n809_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1339gat));
  NOR2_X1   g610(.A1(new_n256_), .A2(new_n495_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n711_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n623_), .A2(new_n625_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n536_), .A2(new_n538_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n533_), .A2(G229gat), .A3(G233gat), .A4(new_n518_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n528_), .A2(new_n518_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n503_), .B1(new_n818_), .B2(new_n519_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT114), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n820_), .A2(KEYINPUT114), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n816_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n815_), .A2(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n592_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(KEYINPUT55), .A4(new_n595_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n607_), .B(new_n604_), .C1(new_n616_), .C2(new_n542_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n594_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT113), .B1(new_n608_), .B2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n828_), .A2(KEYINPUT112), .A3(new_n594_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n827_), .A2(new_n831_), .A3(new_n833_), .A4(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n609_), .A2(new_n614_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n622_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT56), .B(new_n622_), .C1(new_n835_), .C2(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n539_), .A2(new_n625_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT110), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT110), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n539_), .A2(new_n846_), .A3(new_n625_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n824_), .B1(new_n843_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n814_), .B1(new_n849_), .B2(new_n682_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n823_), .A2(new_n625_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n842_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n828_), .A2(KEYINPUT112), .A3(new_n594_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT112), .B1(new_n828_), .B2(new_n594_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n855_), .A2(new_n837_), .A3(new_n833_), .A4(new_n827_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT56), .B1(new_n856_), .B2(new_n622_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n851_), .B1(new_n852_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n843_), .A2(KEYINPUT58), .A3(new_n851_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n661_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n845_), .A2(new_n847_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n864_));
  OAI211_X1 g663(.A(KEYINPUT57), .B(new_n657_), .C1(new_n864_), .C2(new_n824_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n850_), .A2(new_n862_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n850_), .A2(new_n862_), .A3(new_n865_), .A4(KEYINPUT115), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n676_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n661_), .A2(new_n755_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n630_), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n661_), .A2(new_n629_), .A3(KEYINPUT54), .A4(new_n755_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n813_), .B1(new_n870_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G113gat), .B1(new_n877_), .B2(new_n539_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n870_), .A2(new_n876_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n813_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT59), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n866_), .A2(new_n676_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n880_), .B(new_n883_), .C1(new_n884_), .C2(new_n875_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n540_), .A2(KEYINPUT116), .ZN(new_n888_));
  MUX2_X1   g687(.A(KEYINPUT116), .B(new_n888_), .S(G113gat), .Z(new_n889_));
  AOI21_X1  g688(.A(new_n878_), .B1(new_n887_), .B2(new_n889_), .ZN(G1340gat));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n634_), .A2(new_n891_), .ZN(new_n892_));
  MUX2_X1   g691(.A(new_n892_), .B(new_n891_), .S(G120gat), .Z(new_n893_));
  NOR2_X1   g692(.A1(new_n881_), .A2(new_n893_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT117), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n634_), .B(new_n885_), .C1(new_n877_), .C2(new_n883_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(KEYINPUT118), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(KEYINPUT118), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G120gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n895_), .B1(new_n897_), .B2(new_n899_), .ZN(G1341gat));
  OAI211_X1 g699(.A(new_n675_), .B(new_n885_), .C1(new_n877_), .C2(new_n883_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G127gat), .ZN(new_n902_));
  INV_X1    g701(.A(G127gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n877_), .A2(new_n903_), .A3(new_n675_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT119), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n902_), .A2(new_n907_), .A3(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1342gat));
  OAI21_X1  g708(.A(G134gat), .B1(new_n886_), .B2(new_n705_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n657_), .A2(G134gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n881_), .B2(new_n911_), .ZN(G1343gat));
  NOR4_X1   g711(.A1(new_n257_), .A2(new_n498_), .A3(new_n473_), .A4(new_n495_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n879_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT120), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n914_), .A2(KEYINPUT120), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n539_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(G141gat), .ZN(new_n919_));
  INV_X1    g718(.A(G141gat), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n920_), .B(new_n539_), .C1(new_n916_), .C2(new_n917_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1344gat));
  OAI21_X1  g721(.A(new_n634_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT121), .B(G148gat), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n634_), .B(new_n924_), .C1(new_n916_), .C2(new_n917_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1345gat));
  OAI21_X1  g727(.A(new_n675_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT61), .B(G155gat), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n930_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n675_), .B(new_n932_), .C1(new_n916_), .C2(new_n917_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1346gat));
  AND2_X1   g733(.A1(new_n879_), .A2(new_n913_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n705_), .B1(new_n937_), .B2(new_n915_), .ZN(new_n938_));
  INV_X1    g737(.A(G162gat), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n916_), .A2(new_n917_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n682_), .A2(new_n939_), .ZN(new_n941_));
  OAI22_X1  g740(.A1(new_n938_), .A2(new_n939_), .B1(new_n940_), .B2(new_n941_), .ZN(G1347gat));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n884_), .A2(new_n875_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n712_), .A2(new_n498_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n477_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n540_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n943_), .B1(new_n949_), .B2(new_n202_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n949_), .A2(new_n337_), .A3(new_n227_), .ZN(new_n951_));
  OAI211_X1 g750(.A(KEYINPUT62), .B(G169gat), .C1(new_n948_), .C2(new_n540_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n950_), .A2(new_n951_), .A3(new_n952_), .ZN(G1348gat));
  NOR3_X1   g752(.A1(new_n944_), .A2(new_n477_), .A3(new_n946_), .ZN(new_n954_));
  AOI21_X1  g753(.A(G176gat), .B1(new_n954_), .B2(new_n634_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n477_), .B1(new_n870_), .B2(new_n876_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n635_), .A2(new_n203_), .A3(new_n946_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n955_), .B1(new_n956_), .B2(new_n957_), .ZN(G1349gat));
  NAND4_X1  g757(.A1(new_n956_), .A2(new_n498_), .A3(new_n712_), .A4(new_n675_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(new_n342_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n676_), .A2(new_n214_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n945_), .A2(new_n947_), .A3(new_n961_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(KEYINPUT122), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n954_), .A2(new_n964_), .A3(new_n961_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n960_), .A2(new_n963_), .A3(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(KEYINPUT123), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n968_));
  NAND4_X1  g767(.A1(new_n960_), .A2(new_n963_), .A3(new_n968_), .A4(new_n965_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n967_), .A2(new_n969_), .ZN(G1350gat));
  NAND4_X1  g769(.A1(new_n954_), .A2(new_n361_), .A3(new_n362_), .A4(new_n682_), .ZN(new_n971_));
  OAI21_X1  g770(.A(G190gat), .B1(new_n948_), .B2(new_n705_), .ZN(new_n972_));
  AND2_X1   g771(.A1(new_n972_), .A2(KEYINPUT124), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n972_), .A2(KEYINPUT124), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n971_), .B1(new_n973_), .B2(new_n974_), .ZN(G1351gat));
  NAND4_X1  g774(.A1(new_n498_), .A2(new_n495_), .A3(new_n477_), .A4(new_n256_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n976_), .B1(new_n870_), .B2(new_n876_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n977_), .A2(new_n539_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g778(.A1(new_n977_), .A2(new_n634_), .ZN(new_n980_));
  XNOR2_X1  g779(.A(new_n980_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g780(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n982_));
  OAI21_X1  g781(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n983_));
  INV_X1    g782(.A(new_n983_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n984_), .A2(new_n982_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n675_), .A2(new_n986_), .ZN(new_n987_));
  XOR2_X1   g786(.A(new_n987_), .B(KEYINPUT125), .Z(new_n988_));
  NAND2_X1  g787(.A1(new_n977_), .A2(new_n988_), .ZN(new_n989_));
  MUX2_X1   g788(.A(new_n982_), .B(new_n985_), .S(new_n989_), .Z(G1354gat));
  AOI21_X1  g789(.A(G218gat), .B1(new_n977_), .B2(new_n682_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n661_), .A2(G218gat), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n992_), .B(KEYINPUT127), .ZN(new_n993_));
  AOI21_X1  g792(.A(new_n991_), .B1(new_n977_), .B2(new_n993_), .ZN(G1355gat));
endmodule


