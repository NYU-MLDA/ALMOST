//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  OR2_X1    g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  OR3_X1    g006(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n204_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT8), .B1(new_n204_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OAI221_X1 g013(.A(new_n204_), .B1(new_n212_), .B2(KEYINPUT8), .C1(new_n207_), .C2(new_n210_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n207_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT10), .B(G99gat), .Z(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(KEYINPUT9), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(KEYINPUT9), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n221_), .A2(G85gat), .A3(G92gat), .A4(new_n222_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n202_), .A2(new_n220_), .A3(KEYINPUT9), .A4(new_n203_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n216_), .A2(new_n219_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n214_), .A2(new_n215_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n227_));
  AND2_X1   g026(.A1(G71gat), .A2(G78gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G71gat), .A2(G78gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n227_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G57gat), .B(G64gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n228_), .A2(new_n229_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(KEYINPUT11), .ZN(new_n235_));
  INV_X1    g034(.A(G71gat), .ZN(new_n236_));
  INV_X1    g035(.A(G78gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G71gat), .A2(G78gat), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n238_), .A2(new_n233_), .A3(KEYINPUT11), .A4(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n232_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(KEYINPUT11), .A3(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT67), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n244_), .A2(new_n240_), .A3(new_n231_), .A4(new_n230_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n242_), .A2(KEYINPUT68), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT68), .B1(new_n242_), .B2(new_n245_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n226_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT12), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G230gat), .A2(G233gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT64), .Z(new_n252_));
  AND3_X1   g051(.A1(new_n214_), .A2(new_n215_), .A3(new_n225_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n245_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n242_), .A2(KEYINPUT68), .A3(new_n245_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n226_), .A2(KEYINPUT12), .A3(new_n245_), .A4(new_n242_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n250_), .A2(new_n252_), .A3(new_n258_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n248_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n252_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G120gat), .B(G148gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT5), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G176gat), .ZN(new_n266_));
  INV_X1    g065(.A(G204gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n260_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT69), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n260_), .A2(new_n263_), .A3(new_n272_), .A4(new_n269_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n269_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT70), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(new_n279_), .A3(new_n276_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(KEYINPUT13), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT13), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n283_));
  AOI211_X1 g082(.A(KEYINPUT70), .B(new_n275_), .C1(new_n271_), .C2(new_n273_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G113gat), .B(G141gat), .ZN(new_n287_));
  INV_X1    g086(.A(G169gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(G197gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G1gat), .ZN(new_n292_));
  INV_X1    g091(.A(G8gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT14), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT75), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n297_), .B(KEYINPUT14), .C1(new_n292_), .C2(new_n293_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n295_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n299_), .A2(new_n300_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G50gat), .ZN(new_n304_));
  INV_X1    g103(.A(G29gat), .ZN(new_n305_));
  INV_X1    g104(.A(G36gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G43gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G29gat), .A2(G36gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n308_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n304_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G29gat), .B(G36gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G43gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(G50gat), .A3(new_n310_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n303_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n317_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(KEYINPUT81), .A3(new_n320_), .ZN(new_n321_));
  OR3_X1    g120(.A1(new_n303_), .A2(new_n318_), .A3(KEYINPUT81), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G229gat), .A2(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n321_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n303_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT15), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n311_), .A2(new_n304_), .A3(new_n312_), .ZN(new_n328_));
  AOI21_X1  g127(.A(G50gat), .B1(new_n315_), .B2(new_n310_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n313_), .A2(KEYINPUT15), .A3(new_n316_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(new_n323_), .A3(new_n319_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n325_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n291_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  AOI211_X1 g136(.A(KEYINPUT82), .B(new_n290_), .C1(new_n325_), .C2(new_n334_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n286_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G120gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G127gat), .B(G134gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G113gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n342_), .A2(G113gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n341_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n345_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(G120gat), .A3(new_n343_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350_));
  INV_X1    g149(.A(G183gat), .ZN(new_n351_));
  INV_X1    g150(.A(G190gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT24), .ZN(new_n355_));
  INV_X1    g154(.A(G176gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n288_), .A3(new_n356_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n353_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT83), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT25), .B1(new_n359_), .B2(new_n351_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT26), .B1(new_n361_), .B2(new_n352_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT83), .A3(G183gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT26), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n360_), .A2(new_n362_), .A3(new_n364_), .A4(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT85), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n370_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n368_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n358_), .A2(new_n367_), .A3(new_n371_), .A4(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n353_), .B(new_n354_), .C1(G183gat), .C2(G190gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G169gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n349_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G15gat), .B(G43gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT31), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n381_), .B(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G71gat), .B(G99gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT30), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  XOR2_X1   g187(.A(new_n384_), .B(new_n388_), .Z(new_n389_));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n390_), .B(KEYINPUT18), .Z(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G64gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n390_), .B(KEYINPUT18), .ZN(new_n393_));
  INV_X1    g192(.A(G64gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n392_), .A2(new_n395_), .A3(G92gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(G92gat), .B1(new_n392_), .B2(new_n395_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT19), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT92), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n401_), .B(KEYINPUT19), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT92), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n375_), .A2(new_n379_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G211gat), .B(G218gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT88), .B1(new_n267_), .B2(G197gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(KEYINPUT21), .A3(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G197gat), .B(G204gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n414_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n416_), .A2(KEYINPUT21), .A3(new_n411_), .A4(new_n412_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n411_), .A2(KEYINPUT21), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n409_), .B1(new_n410_), .B2(new_n419_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT25), .B(G183gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT26), .B(G190gat), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n422_), .A2(new_n423_), .B1(new_n372_), .B2(new_n368_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n358_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n379_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n408_), .B1(new_n420_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n421_), .A2(new_n380_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n424_), .A2(new_n358_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n409_), .B1(new_n419_), .B2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n431_), .A3(new_n403_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n398_), .B1(new_n428_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n419_), .A2(new_n379_), .A3(new_n375_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n427_), .A2(KEYINPUT20), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n408_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n396_), .A2(new_n397_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n432_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n434_), .A2(new_n435_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT27), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n428_), .A2(new_n433_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(KEYINPUT93), .A3(new_n440_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT98), .B1(new_n444_), .B2(new_n440_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT98), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n441_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT27), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n426_), .A2(KEYINPUT96), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT96), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n430_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n419_), .A3(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n429_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT97), .B1(new_n454_), .B2(KEYINPUT20), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n405_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n437_), .A2(new_n438_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n440_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n446_), .B1(new_n450_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G155gat), .A2(G162gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT86), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G141gat), .A2(G148gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT3), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(KEYINPUT87), .A2(KEYINPUT2), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G141gat), .A2(G148gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(KEYINPUT87), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n471_), .B1(new_n472_), .B2(new_n469_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n464_), .B(new_n465_), .C1(new_n468_), .C2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n466_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT86), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n463_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n465_), .B(KEYINPUT1), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n470_), .B(new_n475_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n349_), .A2(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n346_), .A2(new_n348_), .A3(new_n474_), .A4(new_n479_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(KEYINPUT4), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT4), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n349_), .A2(new_n480_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G225gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G57gat), .B(G85gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n488_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n489_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n487_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n494_), .B1(new_n499_), .B2(new_n496_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G78gat), .B(G106gat), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n419_), .B1(new_n480_), .B2(KEYINPUT29), .ZN(new_n505_));
  OAI211_X1 g304(.A(G228gat), .B(G233gat), .C1(new_n419_), .C2(KEYINPUT89), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n505_), .A2(new_n506_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n504_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n480_), .A2(KEYINPUT29), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT28), .B(G22gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(new_n304_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n513_), .B(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n505_), .A2(new_n506_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n507_), .A3(new_n503_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n512_), .A2(new_n516_), .B1(new_n518_), .B2(new_n510_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n510_), .A2(new_n518_), .A3(KEYINPUT90), .A4(new_n516_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n502_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n462_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n503_), .B1(new_n517_), .B2(new_n507_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n516_), .B1(new_n524_), .B2(KEYINPUT90), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n510_), .A2(new_n518_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n520_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n442_), .A2(new_n445_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n481_), .A2(new_n488_), .A3(new_n482_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n495_), .B(new_n530_), .C1(new_n486_), .C2(new_n488_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT33), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT95), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n494_), .B(new_n533_), .C1(new_n499_), .C2(new_n496_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n500_), .A2(KEYINPUT95), .A3(new_n532_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n529_), .A2(new_n531_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n440_), .A2(KEYINPUT32), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n444_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n454_), .A2(KEYINPUT20), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(new_n429_), .A3(new_n455_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n459_), .B1(new_n542_), .B2(new_n405_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n501_), .B(new_n538_), .C1(new_n543_), .C2(new_n537_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n528_), .B1(new_n536_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n389_), .B1(new_n523_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n462_), .A2(KEYINPUT99), .ZN(new_n547_));
  INV_X1    g346(.A(new_n528_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT99), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n549_), .B(new_n446_), .C1(new_n450_), .C2(new_n461_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n389_), .A2(new_n501_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n547_), .A2(new_n548_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n546_), .A2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n340_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n256_), .A2(new_n257_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT79), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n303_), .B(new_n561_), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n560_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n563_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n562_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n254_), .B(KEYINPUT76), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n573_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n574_), .A2(new_n568_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT35), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n332_), .A2(new_n226_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT72), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n253_), .A2(new_n318_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n588_), .A2(KEYINPUT71), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT71), .ZN(new_n590_));
  AND4_X1   g389(.A1(new_n580_), .A2(new_n586_), .A3(new_n589_), .A4(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n585_), .A2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n586_), .A2(new_n580_), .A3(new_n589_), .A4(new_n590_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT73), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(G134gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(G162gat), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(G162gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n598_), .B(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n602_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT74), .ZN(new_n610_));
  INV_X1    g409(.A(new_n594_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n593_), .B1(new_n584_), .B2(new_n582_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n592_), .A2(KEYINPUT74), .A3(new_n594_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n613_), .A2(new_n601_), .A3(new_n605_), .A4(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n602_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n578_), .B(new_n609_), .C1(new_n608_), .C2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n554_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT100), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n619_), .A2(new_n292_), .A3(new_n501_), .A4(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n620_), .A2(KEYINPUT100), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n617_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(new_n578_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n554_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n501_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT101), .B1(new_n629_), .B2(G1gat), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(KEYINPUT101), .A3(G1gat), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n624_), .B1(new_n630_), .B2(new_n631_), .ZN(G1324gat));
  NAND2_X1  g431(.A1(new_n547_), .A2(new_n550_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n628_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(KEYINPUT102), .A2(KEYINPUT39), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(G8gat), .A3(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(KEYINPUT102), .A2(KEYINPUT39), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n619_), .A2(new_n293_), .A3(new_n633_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n637_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n634_), .A2(G8gat), .A3(new_n635_), .A4(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n389_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n619_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n628_), .B2(new_n646_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(KEYINPUT41), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(KEYINPUT41), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n647_), .B1(new_n649_), .B2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n619_), .A2(new_n652_), .A3(new_n528_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G22gat), .B1(new_n627_), .B2(new_n548_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT42), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(KEYINPUT42), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(G1327gat));
  INV_X1    g456(.A(new_n578_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n617_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n340_), .A2(new_n553_), .A3(new_n659_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(KEYINPUT103), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(KEYINPUT103), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n501_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n305_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n609_), .B1(new_n617_), .B2(new_n608_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n546_), .B2(new_n552_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n340_), .A3(new_n578_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT44), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(G29gat), .A3(new_n501_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n665_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT104), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n679_), .B(new_n665_), .C1(new_n673_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1328gat));
  INV_X1    g480(.A(new_n633_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n671_), .B2(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n675_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n661_), .A2(new_n306_), .A3(new_n633_), .A4(new_n662_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n686_), .A2(new_n687_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n685_), .A2(KEYINPUT46), .A3(new_n688_), .A4(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT46), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n306_), .B1(new_n683_), .B2(new_n675_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n688_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(new_n694_), .ZN(G1329gat));
  NAND4_X1  g494(.A1(new_n672_), .A2(G43gat), .A3(new_n646_), .A4(new_n675_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n663_), .A2(new_n646_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n308_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g499(.A1(new_n672_), .A2(G50gat), .A3(new_n528_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n663_), .A2(new_n528_), .ZN(new_n702_));
  OAI22_X1  g501(.A1(new_n701_), .A2(new_n676_), .B1(G50gat), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(G1331gat));
  INV_X1    g503(.A(new_n339_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n281_), .B2(new_n285_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n553_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n618_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G57gat), .B1(new_n708_), .B2(new_n501_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n707_), .A2(new_n626_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n501_), .A2(G57gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(G1332gat));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n633_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G64gat), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT105), .B(KEYINPUT48), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n708_), .A2(new_n394_), .A3(new_n633_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT106), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(new_n720_), .A3(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1333gat));
  AOI21_X1  g521(.A(new_n236_), .B1(new_n710_), .B2(new_n646_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT49), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n708_), .A2(new_n236_), .A3(new_n646_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1334gat));
  AOI21_X1  g525(.A(new_n237_), .B1(new_n710_), .B2(new_n528_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT50), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n708_), .A2(new_n237_), .A3(new_n528_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT107), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n728_), .A2(new_n732_), .A3(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1335gat));
  AND2_X1   g533(.A1(new_n707_), .A2(new_n659_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n501_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n706_), .B2(new_n578_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n706_), .A2(new_n737_), .A3(new_n578_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n666_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n668_), .B1(new_n553_), .B2(new_n740_), .ZN(new_n741_));
  AOI211_X1 g540(.A(KEYINPUT43), .B(new_n666_), .C1(new_n546_), .C2(new_n552_), .ZN(new_n742_));
  OAI22_X1  g541(.A1(new_n738_), .A2(new_n739_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n501_), .A2(G85gat), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT109), .Z(new_n746_));
  AOI21_X1  g545(.A(new_n736_), .B1(new_n744_), .B2(new_n746_), .ZN(G1336gat));
  AOI21_X1  g546(.A(G92gat), .B1(new_n735_), .B2(new_n633_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n633_), .A2(G92gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n744_), .B2(new_n749_), .ZN(G1337gat));
  INV_X1    g549(.A(G99gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n744_), .B2(new_n646_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n735_), .A2(new_n217_), .A3(new_n646_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754_));
  OAI22_X1  g553(.A1(new_n752_), .A2(new_n753_), .B1(new_n754_), .B2(KEYINPUT51), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(G1338gat));
  OAI21_X1  g556(.A(KEYINPUT111), .B1(new_n743_), .B2(new_n548_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n286_), .A2(new_n339_), .A3(new_n578_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT108), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n760_), .A2(new_n669_), .A3(new_n761_), .A4(new_n528_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(G106gat), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT52), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n758_), .A2(new_n762_), .A3(new_n765_), .A4(G106gat), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n735_), .A2(new_n218_), .A3(new_n528_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT113), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n769_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n767_), .A2(new_n768_), .A3(new_n771_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1339gat));
  NAND4_X1  g574(.A1(new_n618_), .A2(new_n339_), .A3(new_n281_), .A4(new_n285_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n260_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT114), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n260_), .A2(new_n779_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n260_), .A2(new_n783_), .A3(new_n779_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n250_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n262_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n781_), .A2(new_n782_), .A3(new_n784_), .A4(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n268_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT56), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n335_), .A2(new_n291_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n324_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n323_), .B1(new_n333_), .B2(new_n319_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n790_), .B1(new_n793_), .B2(new_n291_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n787_), .A2(new_n795_), .A3(new_n268_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n789_), .A2(new_n274_), .A3(new_n794_), .A4(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n794_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n788_), .B2(KEYINPUT56), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n801_), .A2(KEYINPUT58), .A3(new_n274_), .A4(new_n796_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n740_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n788_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n787_), .A2(KEYINPUT115), .A3(new_n795_), .A4(new_n268_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n339_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n806_), .A2(new_n789_), .A3(new_n807_), .A4(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n794_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n625_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n803_), .A2(new_n804_), .B1(KEYINPUT57), .B2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n799_), .A2(KEYINPUT117), .A3(new_n740_), .A4(new_n802_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n811_), .B2(KEYINPUT57), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n809_), .A2(new_n810_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT116), .B(new_n816_), .C1(new_n817_), .C2(new_n625_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n812_), .A2(new_n813_), .A3(new_n815_), .A4(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n778_), .B1(new_n819_), .B2(new_n578_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n633_), .A2(new_n528_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(new_n501_), .A3(new_n646_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G113gat), .B1(new_n823_), .B2(new_n705_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n803_), .A2(new_n804_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n811_), .A2(KEYINPUT57), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n813_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n818_), .A2(new_n815_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n578_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n778_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n822_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n826_), .A2(new_n803_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n811_), .A2(KEYINPUT57), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n578_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n830_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n832_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n834_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n705_), .A2(G113gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT118), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n824_), .B1(new_n841_), .B2(new_n843_), .ZN(G1340gat));
  OAI211_X1 g643(.A(new_n286_), .B(new_n840_), .C1(new_n823_), .C2(new_n839_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT60), .B1(new_n286_), .B2(new_n341_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n833_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(G120gat), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n833_), .A2(KEYINPUT60), .A3(new_n846_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1341gat));
  INV_X1    g649(.A(G127gat), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n578_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n834_), .A2(new_n840_), .A3(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT119), .B(new_n851_), .C1(new_n833_), .C2(new_n578_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n820_), .A2(new_n578_), .A3(new_n822_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(G127gat), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n853_), .A2(new_n854_), .A3(new_n857_), .ZN(G1342gat));
  AOI21_X1  g657(.A(G134gat), .B1(new_n823_), .B2(new_n625_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n740_), .A2(G134gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n841_), .B2(new_n860_), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n646_), .A2(new_n548_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n682_), .A2(new_n501_), .A3(new_n862_), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT120), .Z(new_n864_));
  NOR2_X1   g663(.A1(new_n820_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n705_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n286_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT121), .B(G148gat), .Z(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1345gat));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n658_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  AOI21_X1  g672(.A(G162gat), .B1(new_n865_), .B2(new_n625_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n666_), .A2(new_n603_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n865_), .B2(new_n875_), .ZN(G1347gat));
  NAND2_X1  g675(.A1(new_n633_), .A2(new_n551_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n339_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT122), .Z(new_n879_));
  NAND3_X1  g678(.A1(new_n838_), .A2(new_n548_), .A3(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(G169gat), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(KEYINPUT62), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(KEYINPUT62), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n877_), .A2(new_n528_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n838_), .A2(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT22), .B(G169gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n705_), .A2(new_n886_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT123), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n882_), .A2(new_n883_), .B1(new_n885_), .B2(new_n888_), .ZN(G1348gat));
  INV_X1    g688(.A(new_n885_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n356_), .A3(new_n286_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n820_), .A2(new_n528_), .A3(new_n877_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n892_), .A2(new_n286_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n893_), .B2(new_n356_), .ZN(G1349gat));
  INV_X1    g693(.A(new_n422_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n838_), .A2(new_n895_), .A3(new_n658_), .A4(new_n884_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT124), .ZN(new_n897_));
  AOI21_X1  g696(.A(G183gat), .B1(new_n892_), .B2(new_n658_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n885_), .B2(new_n666_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n625_), .A2(new_n423_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n885_), .B2(new_n901_), .ZN(G1351gat));
  NOR2_X1   g701(.A1(new_n820_), .A2(new_n501_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n633_), .A2(new_n862_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(new_n705_), .A3(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g706(.A1(new_n903_), .A2(new_n286_), .A3(new_n905_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n267_), .A2(KEYINPUT125), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1353gat));
  NAND3_X1  g709(.A1(new_n903_), .A2(new_n658_), .A3(new_n905_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT63), .B(G211gat), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n911_), .B2(new_n914_), .ZN(G1354gat));
  XOR2_X1   g714(.A(KEYINPUT126), .B(G218gat), .Z(new_n916_));
  AND2_X1   g715(.A1(new_n740_), .A2(new_n916_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n831_), .A2(new_n502_), .A3(new_n905_), .A4(new_n917_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n820_), .A2(new_n501_), .A3(new_n617_), .A4(new_n904_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n916_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(KEYINPUT127), .B(new_n918_), .C1(new_n919_), .C2(new_n916_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1355gat));
endmodule


