//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(G197gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT88), .B1(new_n204_), .B2(G204gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(G197gat), .ZN(new_n208_));
  OAI211_X1 g007(.A(KEYINPUT21), .B(new_n205_), .C1(new_n206_), .C2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(G197gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n204_), .A2(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n210_), .B(new_n211_), .C1(KEYINPUT88), .C2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT21), .B1(new_n206_), .B2(new_n208_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT89), .B1(new_n216_), .B2(new_n214_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n214_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n212_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT89), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n215_), .A2(new_n217_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223_));
  OR2_X1    g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT77), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT23), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n227_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(KEYINPUT23), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n226_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n236_));
  AND2_X1   g035(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n237_));
  AND2_X1   g036(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n239_));
  OAI22_X1  g038(.A1(new_n236_), .A2(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n223_), .B1(new_n235_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT25), .B(G183gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT26), .B(G190gat), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n246_), .A2(new_n247_), .B1(new_n242_), .B2(new_n241_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n233_), .B1(new_n249_), .B2(new_n227_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n248_), .A2(new_n250_), .A3(KEYINPUT93), .A4(new_n226_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G176gat), .ZN(new_n253_));
  AND2_X1   g052(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n256_), .A2(new_n225_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT94), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n229_), .A2(new_n231_), .A3(new_n227_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n228_), .A2(G183gat), .A3(G190gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(G183gat), .B2(G190gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n225_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT94), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n222_), .B1(new_n252_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n226_), .A2(KEYINPUT76), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT76), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n224_), .A2(new_n269_), .A3(KEYINPUT24), .A4(new_n225_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n248_), .A2(new_n268_), .A3(new_n261_), .A4(new_n270_), .ZN(new_n271_));
  OAI22_X1  g070(.A1(new_n232_), .A2(new_n234_), .B1(G183gat), .B2(G190gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n257_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n215_), .A2(new_n217_), .A3(new_n221_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT20), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n203_), .B1(new_n267_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT95), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n240_), .A2(new_n243_), .A3(new_n270_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(KEYINPUT76), .A2(new_n226_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n279_), .A2(new_n280_), .B1(new_n272_), .B2(new_n257_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n278_), .B1(new_n222_), .B2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n274_), .A2(KEYINPUT95), .A3(new_n275_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(KEYINPUT20), .A3(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n252_), .A2(new_n222_), .A3(new_n266_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n203_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n277_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G8gat), .B(G36gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT97), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT96), .B(KEYINPUT18), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n288_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT98), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT79), .B(G127gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(G113gat), .A2(G120gat), .ZN(new_n301_));
  INV_X1    g100(.A(G134gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G113gat), .A2(G120gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n302_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n300_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n306_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(new_n299_), .A3(new_n304_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n311_));
  INV_X1    g110(.A(G155gat), .ZN(new_n312_));
  INV_X1    g111(.A(G162gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n322_));
  NOR3_X1   g121(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT82), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n321_), .B(new_n322_), .C1(new_n323_), .C2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT83), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT83), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n329_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n328_), .A2(new_n330_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n318_), .B1(new_n326_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n319_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n317_), .B(new_n335_), .ZN(new_n336_));
  AOI211_X1 g135(.A(new_n333_), .B(new_n334_), .C1(new_n336_), .C2(new_n316_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n310_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n328_), .A2(new_n330_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n323_), .A2(new_n324_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n316_), .B(new_n317_), .C1(new_n341_), .C2(new_n325_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n316_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n334_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n319_), .A3(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n342_), .A2(new_n345_), .A3(new_n309_), .A4(new_n307_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n338_), .A2(new_n346_), .A3(KEYINPUT4), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n342_), .A2(new_n345_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n310_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n348_), .A3(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G57gat), .B(G85gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n348_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n338_), .A2(new_n346_), .A3(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n347_), .A2(new_n359_), .A3(new_n351_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n338_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n357_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT33), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n358_), .A2(new_n360_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n294_), .B(new_n277_), .C1(new_n284_), .C2(new_n287_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n288_), .A2(KEYINPUT98), .A3(new_n295_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n298_), .A2(new_n366_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n361_), .A2(KEYINPUT33), .A3(new_n362_), .A4(new_n363_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT100), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT101), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n288_), .A2(KEYINPUT98), .A3(new_n295_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT98), .B1(new_n288_), .B2(new_n295_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n367_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT101), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT100), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n370_), .B(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n366_), .A4(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n361_), .A2(new_n362_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n357_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT103), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT103), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n384_), .A3(new_n357_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n364_), .A3(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n294_), .A2(KEYINPUT32), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n266_), .B1(new_n244_), .B2(new_n235_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n388_), .A2(KEYINPUT102), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(KEYINPUT102), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n222_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n284_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n286_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n267_), .A2(new_n276_), .A3(new_n203_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n387_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n386_), .B(new_n395_), .C1(new_n387_), .C2(new_n288_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n372_), .A2(new_n380_), .A3(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G71gat), .B(G99gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G15gat), .B(G43gat), .Z(new_n401_));
  AND2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n400_), .A2(new_n401_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n274_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n281_), .A2(new_n405_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n400_), .B(new_n401_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n271_), .A2(new_n273_), .A3(new_n405_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n405_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n409_), .A2(new_n413_), .A3(KEYINPUT80), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT31), .ZN(new_n415_));
  INV_X1    g214(.A(new_n310_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT31), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n409_), .A2(new_n413_), .A3(KEYINPUT80), .A4(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n415_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n416_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n423_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(new_n222_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT87), .B(G228gat), .ZN(new_n426_));
  OAI211_X1 g225(.A(G233gat), .B(new_n426_), .C1(new_n222_), .C2(KEYINPUT90), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n275_), .B2(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n431_), .B(new_n426_), .C1(new_n424_), .C2(new_n222_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n433_), .B(KEYINPUT91), .Z(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n428_), .A2(new_n432_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT92), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n428_), .A2(new_n432_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n433_), .ZN(new_n439_));
  XOR2_X1   g238(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(new_n349_), .B2(KEYINPUT29), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n342_), .A2(new_n345_), .A3(new_n423_), .A4(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT86), .B(G50gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT84), .B(G22gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n441_), .A2(new_n443_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n428_), .A2(new_n432_), .A3(new_n450_), .A4(new_n435_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n437_), .A2(new_n439_), .A3(new_n449_), .A4(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n436_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n435_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n454_));
  OAI22_X1  g253(.A1(new_n453_), .A2(new_n454_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n422_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n298_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT27), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n295_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(KEYINPUT27), .A3(new_n367_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n421_), .A2(new_n456_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n452_), .B(new_n455_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n386_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n397_), .A2(new_n457_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469_));
  INV_X1    g268(.A(G1gat), .ZN(new_n470_));
  INV_X1    g269(.A(G8gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G8gat), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n474_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G231gat), .A2(G233gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT73), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n477_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G57gat), .ZN(new_n481_));
  INV_X1    g280(.A(G64gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G57gat), .A2(G64gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G71gat), .B(G78gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT11), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(new_n489_), .A3(new_n484_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n485_), .A2(new_n487_), .A3(KEYINPUT11), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n480_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G127gat), .B(G155gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G211gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT16), .B(G183gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n495_), .B1(KEYINPUT17), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n499_), .B(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n495_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT72), .ZN(new_n507_));
  XOR2_X1   g306(.A(G29gat), .B(G36gat), .Z(new_n508_));
  XNOR2_X1  g307(.A(G43gat), .B(G50gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G43gat), .B(G50gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(G29gat), .B(G36gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT15), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G85gat), .ZN(new_n517_));
  INV_X1    g316(.A(G92gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT8), .B1(new_n521_), .B2(KEYINPUT65), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n523_));
  INV_X1    g322(.A(G99gat), .ZN(new_n524_));
  INV_X1    g323(.A(G106gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n526_), .A2(new_n529_), .A3(new_n530_), .A4(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n521_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n522_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT10), .B(G99gat), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n525_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n519_), .A2(KEYINPUT9), .A3(new_n520_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n520_), .A2(KEYINPUT9), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n529_), .A2(new_n530_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n532_), .B(new_n521_), .C1(KEYINPUT65), .C2(KEYINPUT8), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n534_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n516_), .A2(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n514_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n547_), .A2(new_n548_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n550_), .A2(new_n551_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n507_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G190gat), .B(G218gat), .Z(new_n556_));
  XOR2_X1   g355(.A(G134gat), .B(G162gat), .Z(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT36), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n550_), .A2(new_n551_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(KEYINPUT72), .A3(new_n552_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n560_), .A2(new_n563_), .A3(new_n558_), .A4(new_n552_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT37), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n559_), .B(KEYINPUT71), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(new_n564_), .A3(KEYINPUT37), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n468_), .A2(new_n506_), .A3(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n475_), .A2(new_n476_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n510_), .A2(new_n513_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n514_), .B(KEYINPUT15), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n575_), .B(new_n576_), .C1(new_n577_), .C2(new_n573_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n576_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n477_), .A2(new_n514_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n574_), .B1(new_n476_), .B2(new_n475_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n579_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT75), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G169gat), .B(G197gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT75), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n583_), .A2(new_n584_), .A3(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n589_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n590_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n594_));
  AOI211_X1 g393(.A(KEYINPUT74), .B(KEYINPUT75), .C1(new_n578_), .C2(new_n582_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n593_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT69), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G230gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT64), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n542_), .A2(new_n494_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n493_), .A2(new_n534_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(KEYINPUT12), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n542_), .A2(new_n604_), .A3(new_n494_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n600_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n600_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT66), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(KEYINPUT66), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(G204gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT5), .B(G176gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n609_), .A2(new_n610_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n617_));
  OAI22_X1  g416(.A1(new_n616_), .A2(new_n617_), .B1(KEYINPUT67), .B2(KEYINPUT13), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n609_), .A2(new_n610_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n614_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n609_), .A2(new_n610_), .A3(new_n615_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT67), .B(KEYINPUT13), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n620_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(KEYINPUT68), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(KEYINPUT68), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n598_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n625_), .A2(KEYINPUT68), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(KEYINPUT68), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(KEYINPUT69), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n572_), .A2(new_n597_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n386_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n633_), .A2(G1gat), .A3(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n635_), .A2(KEYINPUT38), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(KEYINPUT38), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n629_), .A2(new_n630_), .A3(new_n597_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT104), .ZN(new_n639_));
  INV_X1    g438(.A(new_n565_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n468_), .A2(new_n506_), .A3(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n642_), .A2(new_n386_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n636_), .B(new_n637_), .C1(new_n470_), .C2(new_n643_), .ZN(G1324gat));
  NAND3_X1  g443(.A1(new_n639_), .A2(new_n463_), .A3(new_n641_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n645_), .A2(new_n646_), .A3(G8gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n645_), .B2(G8gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n463_), .A2(new_n471_), .ZN(new_n649_));
  OAI22_X1  g448(.A1(new_n647_), .A2(new_n648_), .B1(new_n633_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(G1325gat));
  OR3_X1    g451(.A1(new_n633_), .A2(G15gat), .A3(new_n421_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n642_), .A2(new_n422_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(new_n654_), .B2(G15gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(G1326gat));
  NAND3_X1  g456(.A1(new_n639_), .A2(new_n456_), .A3(new_n641_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n658_), .A2(new_n659_), .A3(G22gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n658_), .B2(G22gat), .ZN(new_n661_));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n456_), .A2(new_n662_), .ZN(new_n663_));
  OAI22_X1  g462(.A1(new_n660_), .A2(new_n661_), .B1(new_n633_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(G1327gat));
  NOR2_X1   g465(.A1(new_n468_), .A2(new_n505_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n640_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n638_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n386_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT37), .B1(new_n562_), .B2(new_n564_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n570_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(KEYINPUT43), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n397_), .A2(new_n457_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n464_), .A2(new_n467_), .ZN(new_n676_));
  OAI211_X1 g475(.A(KEYINPUT107), .B(new_n674_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n567_), .B2(new_n570_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n671_), .A2(new_n672_), .A3(KEYINPUT106), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n468_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n673_), .A2(KEYINPUT43), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n468_), .B2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n677_), .A2(new_n682_), .A3(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n639_), .A3(new_n506_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n689_), .A2(G29gat), .A3(new_n386_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n686_), .A2(KEYINPUT44), .A3(new_n639_), .A4(new_n506_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n670_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n691_), .A2(new_n463_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n689_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n463_), .B(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n669_), .A2(new_n694_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n669_), .A2(KEYINPUT45), .A3(new_n694_), .A4(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n693_), .B1(new_n696_), .B2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n687_), .A2(new_n688_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n691_), .A2(new_n463_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G36gat), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n708_), .A2(KEYINPUT46), .A3(new_n702_), .A4(new_n703_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(G1329gat));
  NOR3_X1   g509(.A1(new_n668_), .A2(new_n638_), .A3(new_n421_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n711_), .A2(G43gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n691_), .A2(G43gat), .A3(new_n422_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n706_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT47), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n712_), .B(new_n716_), .C1(new_n706_), .C2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1330gat));
  AOI21_X1  g517(.A(G50gat), .B1(new_n669_), .B2(new_n456_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n691_), .A2(G50gat), .A3(new_n456_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n689_), .ZN(G1331gat));
  NOR2_X1   g520(.A1(new_n626_), .A2(new_n627_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n592_), .A2(new_n596_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n572_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G57gat), .B1(new_n726_), .B2(new_n386_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n632_), .A2(new_n597_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n641_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n634_), .A2(new_n481_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(G1332gat));
  NAND3_X1  g530(.A1(new_n726_), .A2(new_n482_), .A3(new_n699_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n729_), .A2(new_n699_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(G64gat), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT48), .B(new_n482_), .C1(new_n729_), .C2(new_n699_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n726_), .A2(new_n738_), .A3(new_n422_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT49), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n729_), .A2(new_n422_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(G71gat), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT49), .B(new_n738_), .C1(new_n729_), .C2(new_n422_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(G1334gat));
  INV_X1    g543(.A(G78gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n726_), .A2(new_n745_), .A3(new_n456_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n729_), .A2(new_n456_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(G78gat), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT50), .B(new_n745_), .C1(new_n729_), .C2(new_n456_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1335gat));
  NOR3_X1   g550(.A1(new_n668_), .A2(new_n597_), .A3(new_n632_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n386_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n724_), .B(new_n506_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n686_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n634_), .A2(new_n517_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n753_), .B1(new_n757_), .B2(new_n758_), .ZN(G1336gat));
  AOI21_X1  g558(.A(G92gat), .B1(new_n752_), .B2(new_n463_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n698_), .A2(new_n518_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n757_), .B2(new_n761_), .ZN(G1337gat));
  NAND2_X1  g561(.A1(new_n757_), .A2(new_n422_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G99gat), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n728_), .A2(new_n667_), .A3(new_n535_), .A4(new_n640_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n421_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n752_), .A2(KEYINPUT110), .A3(new_n535_), .A4(new_n422_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n764_), .A2(new_n769_), .A3(KEYINPUT111), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT51), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n764_), .A2(new_n769_), .A3(KEYINPUT111), .A4(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n686_), .A2(new_n756_), .A3(new_n456_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(KEYINPUT112), .A2(KEYINPUT52), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(G106gat), .A3(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(KEYINPUT112), .A2(KEYINPUT52), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n752_), .A2(new_n525_), .A3(new_n456_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n778_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n775_), .A2(G106gat), .A3(new_n776_), .A4(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n780_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n779_), .A2(new_n785_), .A3(new_n780_), .A4(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT59), .ZN(new_n789_));
  AND4_X1   g588(.A1(KEYINPUT113), .A2(new_n625_), .A3(new_n724_), .A4(new_n505_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n597_), .B1(new_n618_), .B2(new_n624_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT113), .B1(new_n791_), .B2(new_n505_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n673_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT54), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n616_), .A2(new_n617_), .A3(new_n622_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(KEYINPUT67), .A2(KEYINPUT13), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n724_), .B(new_n505_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n791_), .A2(KEYINPUT113), .A3(new_n505_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n673_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n583_), .A2(new_n589_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n575_), .B1(new_n577_), .B2(new_n573_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n579_), .ZN(new_n808_));
  OR3_X1    g607(.A1(new_n580_), .A2(new_n581_), .A3(new_n579_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n593_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n806_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n603_), .A2(new_n605_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n607_), .A3(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n603_), .A2(new_n600_), .A3(new_n605_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n816_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n606_), .A2(new_n817_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n614_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT56), .B(new_n614_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n616_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n813_), .B1(new_n827_), .B2(new_n597_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n805_), .B1(new_n828_), .B2(new_n640_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n616_), .B(new_n724_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT57), .B(new_n565_), .C1(new_n830_), .C2(new_n813_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n826_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n814_), .A2(new_n607_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n817_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(new_n820_), .A3(new_n819_), .A4(new_n818_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT56), .B1(new_n836_), .B2(new_n614_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n621_), .B(new_n811_), .C1(new_n832_), .C2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n827_), .A2(KEYINPUT58), .A3(new_n811_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n571_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n829_), .A2(new_n831_), .A3(new_n842_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n794_), .A2(new_n804_), .B1(new_n843_), .B2(new_n506_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n463_), .A2(new_n634_), .A3(new_n466_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT115), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n789_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n829_), .A2(new_n831_), .A3(new_n842_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n803_), .B1(new_n802_), .B2(new_n673_), .ZN(new_n850_));
  AOI211_X1 g649(.A(KEYINPUT54), .B(new_n571_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n851_));
  OAI22_X1  g650(.A1(new_n849_), .A2(new_n505_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(KEYINPUT59), .A3(new_n846_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n848_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n788_), .B1(new_n854_), .B2(new_n597_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n844_), .A2(new_n847_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(new_n788_), .A3(new_n597_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT116), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n724_), .B1(new_n848_), .B2(new_n853_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n860_), .B(new_n857_), .C1(new_n861_), .C2(new_n788_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(G1340gat));
  NOR2_X1   g662(.A1(new_n722_), .A2(G120gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n856_), .B1(KEYINPUT60), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n632_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n854_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(KEYINPUT60), .B2(new_n865_), .ZN(G1341gat));
  AOI21_X1  g668(.A(G127gat), .B1(new_n856_), .B2(new_n505_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n870_), .A2(KEYINPUT117), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(KEYINPUT117), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n505_), .A2(G127gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT118), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n871_), .A2(new_n872_), .B1(new_n854_), .B2(new_n874_), .ZN(G1342gat));
  AOI21_X1  g674(.A(G134gat), .B1(new_n856_), .B2(new_n640_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n571_), .A2(G134gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT119), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n854_), .B2(new_n878_), .ZN(G1343gat));
  NAND4_X1  g678(.A1(new_n698_), .A2(new_n386_), .A3(new_n456_), .A4(new_n421_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT120), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n844_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n597_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n866_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n505_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  AOI21_X1  g688(.A(G162gat), .B1(new_n882_), .B2(new_n640_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n891_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n681_), .A2(new_n313_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n892_), .A2(new_n893_), .B1(new_n882_), .B2(new_n894_), .ZN(G1347gat));
  NOR4_X1   g694(.A1(new_n844_), .A2(new_n386_), .A3(new_n466_), .A4(new_n698_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n597_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n897_), .A2(G169gat), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n897_), .B2(G169gat), .ZN(new_n900_));
  INV_X1    g699(.A(new_n896_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n597_), .B1(new_n255_), .B2(new_n254_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT123), .ZN(new_n903_));
  OAI22_X1  g702(.A1(new_n899_), .A2(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(G1348gat));
  AOI21_X1  g703(.A(G176gat), .B1(new_n896_), .B2(new_n723_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n896_), .A2(G176gat), .A3(new_n866_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT124), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n896_), .A2(new_n908_), .A3(G176gat), .A4(new_n866_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n905_), .B1(new_n907_), .B2(new_n909_), .ZN(G1349gat));
  NAND2_X1  g709(.A1(new_n896_), .A2(new_n505_), .ZN(new_n911_));
  MUX2_X1   g710(.A(new_n246_), .B(G183gat), .S(new_n911_), .Z(G1350gat));
  OAI21_X1  g711(.A(G190gat), .B1(new_n901_), .B2(new_n673_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n640_), .A2(new_n247_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT125), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n901_), .B2(new_n915_), .ZN(G1351gat));
  NOR4_X1   g715(.A1(new_n844_), .A2(new_n386_), .A3(new_n465_), .A4(new_n698_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n597_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n866_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g720(.A(new_n506_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n922_), .A2(new_n923_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n917_), .A2(new_n925_), .A3(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n927_), .B(new_n928_), .Z(G1354gat));
  AOI21_X1  g728(.A(G218gat), .B1(new_n917_), .B2(new_n640_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n571_), .A2(G218gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n917_), .B2(new_n931_), .ZN(G1355gat));
endmodule


