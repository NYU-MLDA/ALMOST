//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_;
  XNOR2_X1  g000(.A(KEYINPUT10), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT64), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G85gat), .B(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n206_), .A2(KEYINPUT65), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT9), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n210_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT6), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n205_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT68), .ZN(new_n219_));
  INV_X1    g018(.A(G99gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(new_n204_), .A3(KEYINPUT66), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT7), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n223_), .A2(new_n220_), .A3(new_n204_), .A4(KEYINPUT66), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n217_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n207_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT8), .ZN(new_n227_));
  INV_X1    g026(.A(new_n217_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n215_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n219_), .A2(new_n227_), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G29gat), .B(G36gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G43gat), .B(G50gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT15), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G232gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT34), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(KEYINPUT35), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n226_), .A2(KEYINPUT8), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n226_), .A2(KEYINPUT8), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n241_), .A2(new_n242_), .B1(new_n215_), .B2(new_n229_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n240_), .B1(new_n243_), .B2(new_n235_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n237_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n239_), .A2(KEYINPUT35), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n246_), .B(KEYINPUT70), .Z(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n237_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G190gat), .B(G218gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G134gat), .B(G162gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT36), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT73), .B1(new_n251_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT73), .ZN(new_n261_));
  AOI211_X1 g060(.A(new_n261_), .B(new_n258_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n256_), .B(new_n257_), .ZN(new_n263_));
  OAI22_X1  g062(.A1(new_n260_), .A2(new_n262_), .B1(new_n251_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT37), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n251_), .A2(new_n263_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n250_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n247_), .B1(new_n237_), .B2(new_n244_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n259_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n261_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n251_), .A2(KEYINPUT73), .A3(new_n259_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n268_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n265_), .A2(new_n266_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n267_), .A2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G127gat), .B(G155gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT16), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G183gat), .B(G211gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT17), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT78), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n283_), .B2(new_n282_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G57gat), .B(G64gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n290_));
  XOR2_X1   g089(.A(G71gat), .B(G78gat), .Z(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n290_), .A2(new_n291_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(KEYINPUT77), .Z(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(KEYINPUT75), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(KEYINPUT75), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G15gat), .B(G22gat), .ZN(new_n302_));
  INV_X1    g101(.A(G1gat), .ZN(new_n303_));
  INV_X1    g102(.A(G8gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT14), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n299_), .A2(new_n305_), .A3(new_n302_), .A4(new_n300_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT76), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G231gat), .A2(G233gat), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n311_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n297_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n297_), .A3(new_n313_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n288_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n286_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n318_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT79), .B1(new_n317_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n287_), .B1(new_n318_), .B2(new_n314_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n315_), .A2(new_n286_), .A3(new_n316_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT79), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT80), .B1(new_n278_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n227_), .A2(new_n218_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT67), .B1(new_n328_), .B2(new_n296_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n296_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n331_));
  INV_X1    g130(.A(new_n296_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n243_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n329_), .A2(new_n330_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT12), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n296_), .A2(KEYINPUT12), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n330_), .A2(new_n338_), .B1(new_n232_), .B2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n243_), .B2(new_n332_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G120gat), .B(G148gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(G176gat), .B(G204gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n337_), .A2(new_n343_), .A3(new_n349_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT13), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(KEYINPUT13), .A3(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n326_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n359_), .A2(new_n267_), .A3(new_n360_), .A4(new_n277_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n327_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT81), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT18), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT99), .ZN(new_n370_));
  INV_X1    g169(.A(G197gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT93), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT93), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G197gat), .ZN(new_n374_));
  INV_X1    g173(.A(G204gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT21), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(G197gat), .B2(G204gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT94), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n381_), .A3(new_n378_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G211gat), .B(G218gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G197gat), .A2(G204gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT93), .B(G197gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n375_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n385_), .B1(new_n389_), .B2(new_n377_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n389_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n384_), .A2(new_n377_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n383_), .A2(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT26), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT26), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G190gat), .ZN(new_n397_));
  INV_X1    g196(.A(G183gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT25), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT25), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G183gat), .ZN(new_n401_));
  AND4_X1   g200(.A1(new_n395_), .A2(new_n397_), .A3(new_n399_), .A4(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT24), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT24), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n407_), .B2(new_n403_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT23), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT23), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(G183gat), .A3(G190gat), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n402_), .A2(new_n408_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n411_), .A2(KEYINPUT85), .A3(G183gat), .A4(G190gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n410_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT86), .B(G176gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT22), .B(G169gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT98), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n406_), .B(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n414_), .B1(new_n422_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n370_), .B1(new_n393_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n391_), .A2(new_n392_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n376_), .A2(new_n381_), .A3(new_n378_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n381_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n375_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n377_), .B1(new_n435_), .B2(new_n386_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n384_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n431_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n414_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n416_), .A2(new_n417_), .B1(KEYINPUT23), .B2(new_n409_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n425_), .B(new_n427_), .C1(new_n440_), .C2(new_n420_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n442_), .A3(KEYINPUT99), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n430_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT25), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n400_), .A2(KEYINPUT84), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(G183gat), .ZN(new_n448_));
  OR3_X1    g247(.A1(new_n400_), .A2(KEYINPUT83), .A3(G183gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT26), .B(G190gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n399_), .A2(KEYINPUT83), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .A4(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n408_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n419_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n406_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n410_), .A2(new_n412_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(new_n421_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n423_), .A2(new_n424_), .A3(KEYINPUT87), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT87), .B1(new_n423_), .B2(new_n424_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT20), .B1(new_n438_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT97), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n436_), .B(new_n384_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n464_), .A2(new_n431_), .A3(new_n460_), .A4(new_n454_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT97), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(KEYINPUT20), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n444_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G226gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT19), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n461_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT20), .B1(new_n472_), .B2(new_n393_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n470_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n369_), .B1(new_n471_), .B2(new_n477_), .ZN(new_n478_));
  AOI211_X1 g277(.A(new_n368_), .B(new_n476_), .C1(new_n468_), .C2(new_n470_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n364_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n464_), .A2(KEYINPUT96), .A3(new_n431_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT96), .B1(new_n464_), .B2(new_n431_), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n482_), .A2(new_n483_), .A3(new_n442_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n470_), .B1(new_n484_), .B2(new_n473_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n444_), .A2(new_n463_), .A3(new_n474_), .A4(new_n467_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n369_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n471_), .A2(new_n369_), .A3(new_n477_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT27), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n480_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G141gat), .A2(G148gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT2), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT2), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n491_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  OAI22_X1  g295(.A1(KEYINPUT91), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(G141gat), .A2(G148gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n494_), .A2(new_n496_), .A3(new_n497_), .A4(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G155gat), .B(G162gat), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT1), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(G141gat), .B(G148gat), .Z(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT29), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G228gat), .A2(G233gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n438_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT96), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n438_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n516_), .B2(new_n481_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n512_), .B1(new_n517_), .B2(new_n511_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G78gat), .B(G106gat), .Z(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OR3_X1    g319(.A1(new_n509_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT28), .B1(new_n509_), .B2(KEYINPUT29), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G22gat), .B(G50gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n519_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(new_n512_), .C1(new_n517_), .C2(new_n511_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n520_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n525_), .B1(new_n520_), .B2(new_n527_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n490_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G71gat), .B(G99gat), .ZN(new_n533_));
  INV_X1    g332(.A(G43gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT30), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G227gat), .A2(G233gat), .ZN(new_n537_));
  INV_X1    g336(.A(G15gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n536_), .B(new_n539_), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n472_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n536_), .B(new_n539_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n461_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(KEYINPUT90), .A3(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT31), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT31), .ZN(new_n546_));
  INV_X1    g345(.A(G113gat), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(G120gat), .ZN(new_n548_));
  INV_X1    g347(.A(G120gat), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(G113gat), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT88), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(G113gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(G120gat), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G127gat), .B(G134gat), .Z(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT89), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G127gat), .B(G134gat), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n554_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n551_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n559_), .B1(KEYINPUT89), .B2(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n545_), .A2(new_n546_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G1gat), .B(G29gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT103), .B(G85gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT0), .B(G57gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G225gat), .A2(G233gat), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n561_), .A2(new_n562_), .A3(new_n560_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n556_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT89), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n557_), .A2(new_n558_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n509_), .A3(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n565_), .A2(new_n508_), .A3(new_n503_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT4), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT101), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT101), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n581_), .A2(new_n585_), .A3(KEYINPUT4), .A4(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT4), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n579_), .A2(new_n509_), .A3(new_n588_), .A4(new_n580_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT102), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n576_), .B1(new_n587_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n576_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n575_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n566_), .A2(KEYINPUT102), .A3(new_n588_), .A4(new_n509_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT102), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n589_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n574_), .B(new_n595_), .C1(new_n600_), .C2(new_n576_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n594_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n532_), .A2(new_n569_), .A3(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n601_), .B(new_n594_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n465_), .A2(new_n466_), .A3(KEYINPUT20), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n466_), .B1(new_n465_), .B2(KEYINPUT20), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n474_), .B1(new_n608_), .B2(new_n444_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n368_), .B1(new_n609_), .B2(new_n476_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT27), .B1(new_n610_), .B2(new_n488_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n479_), .A2(new_n487_), .A3(new_n364_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n605_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n485_), .A2(new_n486_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(KEYINPUT32), .A3(new_n369_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n369_), .A2(KEYINPUT32), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n471_), .A2(new_n616_), .A3(new_n477_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n602_), .A2(new_n615_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n610_), .A2(KEYINPUT100), .A3(new_n488_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OAI211_X1 g421(.A(KEYINPUT33), .B(new_n575_), .C1(new_n591_), .C2(new_n593_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n587_), .A2(new_n590_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n592_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n574_), .B1(new_n625_), .B2(new_n595_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n587_), .A2(new_n576_), .A3(new_n590_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n581_), .A2(new_n592_), .A3(new_n582_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(new_n574_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n627_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n623_), .B1(new_n626_), .B2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n618_), .B1(new_n622_), .B2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n613_), .B1(new_n633_), .B2(new_n530_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n604_), .B1(new_n634_), .B2(new_n569_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n307_), .A2(new_n308_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n636_), .A2(new_n235_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n307_), .A2(new_n235_), .A3(new_n308_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n236_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n639_), .B(new_n641_), .C1(new_n644_), .C2(new_n636_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G113gat), .B(G141gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G169gat), .B(G197gat), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n647_), .B(new_n648_), .Z(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n646_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT82), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n635_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT81), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n327_), .A2(new_n358_), .A3(new_n655_), .A4(new_n361_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n363_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n303_), .A3(new_n602_), .ZN(new_n658_));
  XOR2_X1   g457(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n635_), .A2(KEYINPUT105), .A3(new_n264_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT105), .B1(new_n635_), .B2(new_n264_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n358_), .A2(new_n651_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n317_), .A2(new_n320_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(new_n602_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n660_), .B1(new_n669_), .B2(new_n303_), .ZN(G1324gat));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n490_), .B(new_n667_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n671_), .B1(new_n673_), .B2(new_n304_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n654_), .A2(new_n656_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n490_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(G8gat), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n675_), .A2(KEYINPUT106), .A3(new_n363_), .A4(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n363_), .A2(new_n654_), .A3(new_n656_), .A4(new_n677_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n672_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n674_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1325gat));
  NAND3_X1  g485(.A1(new_n657_), .A2(new_n538_), .A3(new_n569_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n569_), .B(new_n667_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n688_), .B2(G15gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT108), .ZN(G1326gat));
  INV_X1    g491(.A(G22gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n657_), .A2(new_n693_), .A3(new_n531_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n663_), .A2(new_n531_), .A3(new_n667_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G22gat), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(KEYINPUT42), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(KEYINPUT42), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1327gat));
  NOR2_X1   g498(.A1(new_n664_), .A2(new_n359_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n267_), .A2(new_n277_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n569_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n628_), .A2(new_n630_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n594_), .B1(new_n703_), .B2(new_n627_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n704_), .A2(new_n620_), .A3(new_n623_), .A4(new_n621_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n531_), .B1(new_n705_), .B2(new_n618_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n706_), .B2(new_n613_), .ZN(new_n707_));
  AOI211_X1 g506(.A(KEYINPUT43), .B(new_n701_), .C1(new_n707_), .C2(new_n604_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n635_), .B2(new_n278_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n700_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(KEYINPUT44), .B(new_n700_), .C1(new_n708_), .C2(new_n710_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n713_), .A2(G29gat), .A3(new_n602_), .A4(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(G29gat), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n326_), .A2(new_n274_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n357_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n633_), .A2(new_n530_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n613_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n569_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n604_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n653_), .B(new_n718_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n635_), .A2(KEYINPUT109), .A3(new_n653_), .A4(new_n718_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n716_), .B1(new_n727_), .B2(new_n603_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n715_), .A2(new_n728_), .ZN(G1328gat));
  NAND3_X1  g528(.A1(new_n713_), .A2(new_n490_), .A3(new_n714_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G36gat), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n676_), .A2(G36gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n725_), .A2(new_n726_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT110), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n725_), .A2(new_n736_), .A3(new_n726_), .A4(new_n732_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n734_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n735_), .B1(new_n734_), .B2(new_n737_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n731_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n731_), .B(KEYINPUT46), .C1(new_n738_), .C2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1329gat));
  NAND4_X1  g543(.A1(new_n713_), .A2(G43gat), .A3(new_n569_), .A4(new_n714_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n534_), .B1(new_n727_), .B2(new_n702_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g547(.A1(new_n713_), .A2(G50gat), .A3(new_n531_), .A4(new_n714_), .ZN(new_n749_));
  INV_X1    g548(.A(G50gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(new_n727_), .B2(new_n530_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1331gat));
  AND2_X1   g551(.A1(new_n327_), .A2(new_n361_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n357_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n651_), .B1(new_n707_), .B2(new_n604_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n753_), .A2(KEYINPUT111), .A3(new_n357_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n756_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  OR3_X1    g558(.A1(new_n759_), .A2(G57gat), .A3(new_n603_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n358_), .A2(new_n326_), .A3(new_n653_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n663_), .A2(new_n602_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G57gat), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(new_n763_), .ZN(G1332gat));
  OR3_X1    g563(.A1(new_n759_), .A2(G64gat), .A3(new_n676_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n663_), .A2(new_n490_), .A3(new_n761_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G64gat), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(KEYINPUT48), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(KEYINPUT48), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(G1333gat));
  OAI211_X1 g569(.A(new_n569_), .B(new_n761_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(G71gat), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G71gat), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n702_), .A2(G71gat), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n773_), .A2(new_n774_), .B1(new_n759_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT113), .ZN(G1334gat));
  NAND3_X1  g576(.A1(new_n663_), .A2(new_n531_), .A3(new_n761_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G78gat), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(KEYINPUT50), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(KEYINPUT50), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n530_), .A2(G78gat), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT114), .ZN(new_n783_));
  OAI22_X1  g582(.A1(new_n780_), .A2(new_n781_), .B1(new_n759_), .B2(new_n783_), .ZN(G1335gat));
  NOR3_X1   g583(.A1(new_n358_), .A2(new_n359_), .A3(new_n651_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n603_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n717_), .A2(new_n358_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n757_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(new_n212_), .A3(new_n602_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n787_), .A2(new_n790_), .ZN(G1336gat));
  AOI21_X1  g590(.A(G92gat), .B1(new_n789_), .B2(new_n490_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n786_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n490_), .A2(G92gat), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT115), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n792_), .B1(new_n793_), .B2(new_n795_), .ZN(G1337gat));
  NAND4_X1  g595(.A1(new_n757_), .A2(new_n569_), .A3(new_n203_), .A4(new_n788_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT116), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n793_), .A2(new_n569_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(G99gat), .ZN(new_n800_));
  XOR2_X1   g599(.A(new_n800_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g600(.A1(new_n789_), .A2(new_n204_), .A3(new_n531_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n531_), .B(new_n785_), .C1(new_n708_), .C2(new_n710_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n803_), .A2(G106gat), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n803_), .B2(G106gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n802_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g608(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n326_), .A2(new_n653_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n358_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n813_), .B2(new_n278_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n701_), .A2(new_n358_), .A3(new_n812_), .A4(new_n810_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n341_), .A2(KEYINPUT55), .A3(new_n342_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n343_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n341_), .A2(KEYINPUT119), .A3(KEYINPUT55), .A4(new_n342_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n330_), .A2(new_n338_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n232_), .A2(new_n340_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n824_), .A2(new_n329_), .A3(new_n333_), .A4(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n336_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .A4(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n350_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n828_), .A2(KEYINPUT56), .A3(new_n350_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(KEYINPUT120), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n828_), .A2(new_n834_), .A3(KEYINPUT56), .A4(new_n350_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n651_), .A2(new_n352_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n641_), .B(new_n638_), .C1(new_n236_), .C2(new_n309_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n640_), .A2(new_n641_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT121), .A3(new_n650_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n642_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n649_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n838_), .B1(new_n840_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n646_), .A2(new_n650_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n833_), .A2(new_n837_), .B1(new_n353_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n817_), .B1(new_n850_), .B2(new_n274_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n353_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n828_), .A2(KEYINPUT56), .A3(new_n350_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT56), .B1(new_n828_), .B2(new_n350_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n834_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n835_), .A2(new_n836_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n852_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(KEYINPUT57), .A3(new_n264_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n846_), .A2(new_n352_), .A3(new_n848_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n860_), .A2(KEYINPUT58), .B1(new_n277_), .B2(new_n267_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n853_), .A2(new_n854_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n859_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n861_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n851_), .A2(new_n858_), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n816_), .B1(new_n866_), .B2(new_n666_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n702_), .A2(new_n603_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n532_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(new_n547_), .A3(new_n651_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n866_), .A2(new_n326_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n816_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n869_), .A2(KEYINPUT59), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT59), .B1(new_n867_), .B2(new_n869_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n653_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n871_), .B1(new_n878_), .B2(new_n547_), .ZN(G1340gat));
  OAI21_X1  g678(.A(new_n549_), .B1(new_n358_), .B2(KEYINPUT60), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n870_), .B(new_n880_), .C1(KEYINPUT60), .C2(new_n549_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n876_), .A2(new_n877_), .A3(new_n357_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n549_), .ZN(G1341gat));
  INV_X1    g682(.A(G127gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n666_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n876_), .A2(new_n877_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n869_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n857_), .A2(new_n264_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n888_), .A2(new_n817_), .B1(new_n864_), .B2(new_n861_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n665_), .B1(new_n889_), .B2(new_n858_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n359_), .B(new_n887_), .C1(new_n890_), .C2(new_n816_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n884_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n886_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n886_), .A2(new_n892_), .A3(KEYINPUT123), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1342gat));
  INV_X1    g696(.A(G134gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n870_), .A2(new_n898_), .A3(new_n274_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n876_), .A2(new_n877_), .A3(new_n278_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n898_), .ZN(G1343gat));
  NOR4_X1   g700(.A1(new_n569_), .A2(new_n490_), .A3(new_n603_), .A4(new_n530_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n867_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n651_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT124), .B(G141gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1344gat));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n357_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(G148gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1345gat));
  NAND2_X1  g709(.A1(new_n904_), .A2(new_n359_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1346gat));
  INV_X1    g712(.A(G162gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n904_), .A2(new_n914_), .A3(new_n274_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n867_), .A2(new_n701_), .A3(new_n903_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n914_), .ZN(G1347gat));
  NOR3_X1   g716(.A1(new_n702_), .A2(new_n602_), .A3(new_n676_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n531_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n651_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n923_), .A2(new_n924_), .A3(G169gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n923_), .B2(G169gat), .ZN(new_n926_));
  INV_X1    g725(.A(new_n922_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n651_), .A2(new_n424_), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT126), .Z(new_n929_));
  OAI22_X1  g728(.A1(new_n925_), .A2(new_n926_), .B1(new_n927_), .B2(new_n929_), .ZN(G1348gat));
  NAND2_X1  g729(.A1(new_n922_), .A2(new_n357_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n867_), .A2(new_n531_), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n918_), .A2(G176gat), .A3(new_n357_), .ZN(new_n933_));
  AOI22_X1  g732(.A1(new_n931_), .A2(new_n423_), .B1(new_n932_), .B2(new_n933_), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n932_), .A2(new_n359_), .A3(new_n918_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n666_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n935_), .A2(new_n398_), .B1(new_n922_), .B2(new_n936_), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n922_), .A2(new_n450_), .A3(new_n274_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n922_), .A2(new_n278_), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n939_), .A2(KEYINPUT127), .A3(G190gat), .ZN(new_n940_));
  AOI21_X1  g739(.A(KEYINPUT127), .B1(new_n939_), .B2(G190gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n938_), .B1(new_n940_), .B2(new_n941_), .ZN(G1351gat));
  NOR3_X1   g741(.A1(new_n569_), .A2(new_n676_), .A3(new_n605_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n867_), .A2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n651_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n357_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g748(.A1(new_n945_), .A2(new_n665_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  AND2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n950_), .A2(new_n951_), .A3(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n953_), .B1(new_n950_), .B2(new_n951_), .ZN(G1354gat));
  INV_X1    g753(.A(G218gat), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n945_), .A2(new_n955_), .A3(new_n274_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n867_), .A2(new_n701_), .A3(new_n944_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n957_), .B2(new_n955_), .ZN(G1355gat));
endmodule


