//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G113gat), .ZN(new_n203_));
  INV_X1    g002(.A(G120gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G99gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G227gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT30), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n207_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT24), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  MUX2_X1   g013(.A(new_n213_), .B(KEYINPUT24), .S(new_n214_), .Z(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT23), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT79), .B1(new_n219_), .B2(G190gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n218_), .B(new_n220_), .C1(new_n221_), .C2(KEYINPUT79), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n215_), .A2(new_n217_), .A3(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT22), .B(G169gat), .Z(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(G176gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n211_), .A2(new_n212_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT80), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n217_), .A2(KEYINPUT81), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n216_), .A2(KEYINPUT23), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT81), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n227_), .A2(KEYINPUT80), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n223_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G15gat), .B(G43gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n210_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G197gat), .A2(G204gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(KEYINPUT85), .B(G197gat), .Z(new_n244_));
  OAI211_X1 g043(.A(KEYINPUT21), .B(new_n243_), .C1(new_n244_), .C2(G204gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G211gat), .B(G218gat), .ZN(new_n246_));
  INV_X1    g045(.A(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G197gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n245_), .B(new_n246_), .C1(new_n249_), .C2(KEYINPUT21), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n250_), .A2(KEYINPUT86), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(KEYINPUT86), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n246_), .B(KEYINPUT87), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(KEYINPUT21), .A3(new_n249_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G155gat), .B(G162gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT84), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT3), .Z(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT2), .Z(new_n262_));
  OAI21_X1  g061(.A(new_n258_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n264_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n265_));
  OAI221_X1 g064(.A(new_n265_), .B1(G141gat), .B2(G148gat), .C1(KEYINPUT1), .C2(new_n256_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT29), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n255_), .A2(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(G228gat), .A2(G233gat), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(KEYINPUT88), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(KEYINPUT88), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G78gat), .B(G106gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n276_), .B(KEYINPUT89), .Z(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT90), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n272_), .B(new_n277_), .C1(new_n269_), .C2(new_n274_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n267_), .A2(KEYINPUT29), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G22gat), .B(G50gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT28), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n283_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n282_), .B(new_n287_), .C1(new_n280_), .C2(new_n279_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n279_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT91), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT91), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n279_), .A2(new_n291_), .A3(new_n281_), .A4(new_n286_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n288_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G8gat), .B(G36gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(G64gat), .B(G92gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT96), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n299_), .A2(KEYINPUT96), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n221_), .B(KEYINPUT92), .Z(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n218_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n303_), .A2(new_n215_), .A3(new_n233_), .A4(new_n229_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n224_), .B(KEYINPUT93), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n212_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n226_), .B1(new_n217_), .B2(new_n231_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n255_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n255_), .A2(new_n237_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(KEYINPUT20), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT19), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n255_), .A2(new_n309_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n316_), .B(KEYINPUT20), .C1(new_n255_), .C2(new_n237_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n317_), .A2(new_n314_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n300_), .B(new_n301_), .C1(new_n315_), .C2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n314_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n314_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n310_), .A2(KEYINPUT20), .A3(new_n321_), .A4(new_n311_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n320_), .A2(new_n299_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n319_), .A2(new_n324_), .A3(KEYINPUT27), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT27), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n299_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(new_n323_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n205_), .A2(new_n267_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n205_), .A2(new_n267_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n205_), .A2(new_n267_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n205_), .A2(new_n267_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(KEYINPUT4), .A3(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(KEYINPUT4), .B2(new_n337_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n339_), .B2(new_n334_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT0), .B(G57gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(G85gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n340_), .B(new_n344_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n293_), .A2(new_n329_), .A3(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n288_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n323_), .A2(new_n327_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT33), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n332_), .A2(new_n334_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n344_), .B(new_n352_), .C1(new_n339_), .C2(new_n334_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT33), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n349_), .B(new_n354_), .C1(new_n340_), .C2(new_n344_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n348_), .A2(new_n351_), .A3(new_n353_), .A4(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n320_), .A2(new_n322_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n299_), .A2(KEYINPUT32), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n315_), .A2(new_n318_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n345_), .B(new_n359_), .C1(new_n358_), .C2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n347_), .B1(new_n356_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n242_), .B1(new_n346_), .B2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n329_), .A2(new_n347_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n242_), .A2(new_n345_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(KEYINPUT66), .B(G106gat), .Z(new_n368_));
  INV_X1    g167(.A(G99gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT10), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(G99gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT65), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n370_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n368_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT67), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT68), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT9), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(G85gat), .ZN(new_n380_));
  INV_X1    g179(.A(G85gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT68), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G92gat), .ZN(new_n384_));
  INV_X1    g183(.A(G92gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G85gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n381_), .A2(G92gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT9), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G99gat), .A2(G106gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT6), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n384_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT67), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n393_), .B(new_n368_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n377_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT69), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT69), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n377_), .A2(new_n392_), .A3(new_n397_), .A4(new_n394_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n399_));
  OR3_X1    g198(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n391_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n388_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n388_), .A2(KEYINPUT70), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT8), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n401_), .A2(new_n404_), .A3(new_n388_), .A4(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n396_), .A2(new_n398_), .A3(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G57gat), .B(G64gat), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n410_), .A2(KEYINPUT11), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(KEYINPUT11), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G71gat), .B(G78gat), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT72), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT12), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G230gat), .A2(G233gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n419_), .B(KEYINPUT64), .Z(new_n420_));
  OR2_X1    g219(.A1(new_n409_), .A2(new_n415_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT12), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n416_), .A2(KEYINPUT72), .A3(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .A4(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n421_), .A2(new_n425_), .A3(new_n416_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n420_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n409_), .A2(KEYINPUT71), .A3(new_n415_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G120gat), .B(G148gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(new_n247_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT5), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(new_n212_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n430_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT73), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n424_), .A2(new_n429_), .A3(new_n434_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n430_), .A2(KEYINPUT73), .A3(new_n435_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT13), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(KEYINPUT13), .A3(new_n440_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G29gat), .B(G36gat), .ZN(new_n447_));
  INV_X1    g246(.A(G43gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G50gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G15gat), .B(G22gat), .ZN(new_n452_));
  INV_X1    g251(.A(G1gat), .ZN(new_n453_));
  INV_X1    g252(.A(G8gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT14), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G1gat), .B(G8gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n451_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT77), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n451_), .B(KEYINPUT15), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n458_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G229gat), .A2(G233gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(new_n461_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n451_), .A2(KEYINPUT77), .A3(new_n459_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n451_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n467_), .A2(new_n468_), .B1(new_n458_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n466_), .B1(new_n470_), .B2(new_n465_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(G197gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT78), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(new_n211_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n466_), .B(new_n475_), .C1(new_n470_), .C2(new_n465_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n446_), .A2(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n367_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n463_), .A2(new_n409_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n409_), .A2(new_n469_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G232gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT34), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(new_n484_), .A3(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n487_), .A2(new_n488_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n491_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT75), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT74), .B(G134gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G162gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G190gat), .B(G218gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT36), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n492_), .A2(new_n493_), .A3(new_n499_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n495_), .A2(new_n504_), .A3(new_n500_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n502_), .A2(KEYINPUT37), .A3(new_n503_), .A4(new_n505_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G231gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n458_), .B(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n512_), .A2(new_n415_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n415_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT76), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT16), .B(G183gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(G211gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(G127gat), .B(G155gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  OR3_X1    g318(.A1(new_n515_), .A2(KEYINPUT17), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n513_), .A2(new_n514_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n519_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n522_), .B(KEYINPUT17), .C1(new_n515_), .C2(new_n519_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n510_), .A2(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n482_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n453_), .A3(new_n345_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT97), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT38), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n529_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n506_), .A2(new_n524_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n482_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT98), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n482_), .A2(new_n535_), .A3(new_n532_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n345_), .ZN(new_n539_));
  OAI21_X1  g338(.A(G1gat), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n530_), .A2(new_n531_), .A3(new_n540_), .ZN(G1324gat));
  NAND3_X1  g340(.A1(new_n526_), .A2(new_n454_), .A3(new_n329_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT39), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n482_), .A2(new_n329_), .A3(new_n532_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT99), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n544_), .A2(new_n545_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n543_), .B1(new_n548_), .B2(G8gat), .ZN(new_n549_));
  NOR4_X1   g348(.A1(new_n546_), .A2(new_n547_), .A3(KEYINPUT39), .A4(new_n454_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n542_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT40), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(KEYINPUT40), .B(new_n542_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(G1325gat));
  INV_X1    g354(.A(G15gat), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n537_), .B2(new_n241_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT41), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n526_), .A2(new_n556_), .A3(new_n241_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(G1326gat));
  INV_X1    g359(.A(G22gat), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n526_), .A2(new_n561_), .A3(new_n347_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n293_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n563_));
  OR3_X1    g362(.A1(new_n563_), .A2(KEYINPUT100), .A3(new_n561_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT100), .B1(new_n563_), .B2(new_n561_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n564_), .A2(KEYINPUT42), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT42), .B1(new_n564_), .B2(new_n565_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n562_), .B1(new_n566_), .B2(new_n567_), .ZN(G1327gat));
  INV_X1    g367(.A(KEYINPUT43), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n325_), .A2(new_n328_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n539_), .A3(new_n347_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n361_), .A2(new_n356_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n293_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n241_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n366_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n569_), .B(new_n510_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT101), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n574_), .A2(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n508_), .A2(new_n509_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT43), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n367_), .A2(KEYINPUT101), .A3(new_n569_), .A4(new_n510_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n481_), .A3(new_n524_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n583_), .A2(new_n481_), .A3(new_n524_), .A4(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n345_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(G29gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n506_), .A2(new_n524_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT103), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n482_), .A2(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(G29gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n590_), .B1(new_n539_), .B2(new_n594_), .ZN(G1328gat));
  NAND3_X1  g394(.A1(new_n586_), .A2(new_n329_), .A3(new_n588_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(G36gat), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n593_), .A2(G36gat), .A3(new_n570_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT45), .Z(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT46), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n599_), .A3(KEYINPUT46), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1329gat));
  NAND4_X1  g403(.A1(new_n586_), .A2(G43gat), .A3(new_n241_), .A4(new_n588_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n448_), .B1(new_n593_), .B2(new_n242_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g407(.A1(new_n586_), .A2(G50gat), .A3(new_n347_), .A4(new_n588_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n450_), .B1(new_n593_), .B2(new_n293_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT104), .ZN(G1331gat));
  NOR2_X1   g411(.A1(new_n445_), .A2(new_n479_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n579_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n615_), .A2(new_n525_), .ZN(new_n616_));
  AOI21_X1  g415(.A(G57gat), .B1(new_n616_), .B2(new_n345_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n615_), .A2(new_n532_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(G57gat), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(KEYINPUT105), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622_));
  OAI21_X1  g421(.A(G57gat), .B1(new_n539_), .B2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n617_), .B1(new_n621_), .B2(new_n623_), .ZN(G1332gat));
  OAI21_X1  g423(.A(G64gat), .B1(new_n619_), .B2(new_n570_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT106), .Z(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT48), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n625_), .B(KEYINPUT106), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT48), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(G64gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n616_), .A2(new_n631_), .A3(new_n329_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n627_), .A2(new_n630_), .A3(new_n632_), .ZN(G1333gat));
  OAI21_X1  g432(.A(G71gat), .B1(new_n619_), .B2(new_n242_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT107), .Z(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT49), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n634_), .B(KEYINPUT107), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT49), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(G71gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n616_), .A2(new_n640_), .A3(new_n241_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n636_), .A2(new_n639_), .A3(new_n641_), .ZN(G1334gat));
  INV_X1    g441(.A(G78gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n616_), .A2(new_n643_), .A3(new_n347_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G78gat), .B1(new_n619_), .B2(new_n293_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n645_), .A2(KEYINPUT108), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(KEYINPUT108), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n646_), .A2(KEYINPUT50), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT50), .B1(new_n646_), .B2(new_n647_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n644_), .B1(new_n648_), .B2(new_n649_), .ZN(G1335gat));
  AND2_X1   g449(.A1(new_n615_), .A2(new_n592_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G85gat), .B1(new_n651_), .B2(new_n345_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n583_), .A2(new_n524_), .A3(new_n613_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n378_), .A2(G85gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n539_), .B1(new_n382_), .B2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n652_), .B1(new_n653_), .B2(new_n655_), .ZN(G1336gat));
  AOI21_X1  g455(.A(G92gat), .B1(new_n651_), .B2(new_n329_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n653_), .A2(new_n329_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(G92gat), .ZN(G1337gat));
  OAI211_X1 g458(.A(new_n651_), .B(new_n241_), .C1(new_n375_), .C2(new_n374_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT109), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n653_), .A2(new_n241_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G99gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT51), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT51), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(new_n667_), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1338gat));
  NAND3_X1  g468(.A1(new_n651_), .A2(new_n368_), .A3(new_n347_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n583_), .A2(new_n347_), .A3(new_n524_), .A4(new_n613_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT52), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n671_), .A2(new_n672_), .A3(G106gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n671_), .B2(G106gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g475(.A1(KEYINPUT112), .A2(KEYINPUT54), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n477_), .A2(new_n478_), .A3(new_n523_), .A4(new_n520_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n444_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT13), .B1(new_n439_), .B2(new_n440_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(KEYINPUT111), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT111), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n445_), .B2(new_n681_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n580_), .B(new_n678_), .C1(new_n685_), .C2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n684_), .A2(KEYINPUT111), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n445_), .A2(new_n686_), .A3(new_n681_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n510_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n465_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n462_), .A2(new_n464_), .A3(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n695_), .B(new_n476_), .C1(new_n470_), .C2(new_n694_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(new_n478_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(KEYINPUT116), .A3(new_n438_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n438_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT116), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT113), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n422_), .B1(new_n416_), .B2(KEYINPUT72), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT72), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n704_), .B(KEYINPUT12), .C1(new_n409_), .C2(new_n415_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n409_), .A2(new_n415_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n703_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n707_), .B2(new_n420_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(KEYINPUT55), .A3(new_n420_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n418_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(KEYINPUT113), .A3(new_n427_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT55), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n424_), .A2(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n708_), .A2(new_n709_), .A3(new_n711_), .A4(new_n713_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n714_), .A2(KEYINPUT56), .A3(new_n435_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT56), .B1(new_n714_), .B2(new_n435_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n698_), .B(new_n701_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n714_), .A2(new_n435_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT56), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n714_), .A2(KEYINPUT56), .A3(new_n435_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n718_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(new_n701_), .A4(new_n698_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n510_), .A2(new_n719_), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT118), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT57), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n439_), .A2(new_n440_), .A3(new_n697_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n439_), .A2(KEYINPUT115), .A3(new_n440_), .A4(new_n697_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n716_), .A2(KEYINPUT114), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n723_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n714_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n435_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n479_), .A3(new_n438_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n735_), .B1(new_n737_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n730_), .B1(new_n741_), .B2(new_n506_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n506_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n739_), .B1(new_n723_), .B2(new_n736_), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT57), .B(new_n743_), .C1(new_n744_), .C2(new_n735_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n510_), .A2(new_n719_), .A3(new_n726_), .A4(KEYINPUT118), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n729_), .A2(new_n742_), .A3(new_n745_), .A4(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n693_), .B1(new_n747_), .B2(new_n524_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n364_), .A2(new_n345_), .A3(new_n241_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT119), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G113gat), .B1(new_n751_), .B2(new_n479_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT59), .B1(new_n748_), .B2(new_n750_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n693_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n742_), .A2(new_n745_), .A3(new_n727_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n524_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n750_), .A2(KEYINPUT59), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n753_), .A2(KEYINPUT120), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT120), .B1(new_n753_), .B2(new_n759_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n480_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n752_), .B1(new_n762_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g562(.A(new_n204_), .B1(new_n445_), .B2(KEYINPUT60), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n751_), .B(new_n764_), .C1(KEYINPUT60), .C2(new_n204_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n753_), .A2(new_n446_), .A3(new_n759_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n204_), .ZN(G1341gat));
  AOI21_X1  g566(.A(G127gat), .B1(new_n751_), .B2(new_n756_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n760_), .A2(new_n761_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n756_), .A2(G127gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(G1342gat));
  AOI21_X1  g570(.A(G134gat), .B1(new_n751_), .B2(new_n506_), .ZN(new_n772_));
  INV_X1    g571(.A(G134gat), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n760_), .A2(new_n761_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n774_), .B2(new_n510_), .ZN(G1343gat));
  NAND2_X1  g574(.A1(new_n570_), .A2(new_n347_), .ZN(new_n776_));
  NOR4_X1   g575(.A1(new_n748_), .A2(new_n539_), .A3(new_n776_), .A4(new_n241_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n479_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n446_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g580(.A1(new_n777_), .A2(new_n756_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(KEYINPUT61), .B(G155gat), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT121), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n782_), .B(new_n784_), .ZN(G1346gat));
  AOI21_X1  g584(.A(G162gat), .B1(new_n777_), .B2(new_n506_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n510_), .A2(G162gat), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT122), .Z(new_n788_));
  AOI21_X1  g587(.A(new_n786_), .B1(new_n777_), .B2(new_n788_), .ZN(G1347gat));
  AND3_X1   g588(.A1(new_n293_), .A2(new_n329_), .A3(new_n365_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n757_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT123), .B1(new_n791_), .B2(new_n480_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT123), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n757_), .A2(new_n793_), .A3(new_n479_), .A4(new_n790_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(G169gat), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT62), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n791_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n479_), .A3(new_n305_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n792_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n794_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n797_), .A2(new_n799_), .A3(new_n800_), .ZN(G1348gat));
  INV_X1    g600(.A(new_n748_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(new_n790_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n445_), .A2(new_n212_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n803_), .A2(KEYINPUT124), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT124), .B1(new_n803_), .B2(new_n804_), .ZN(new_n806_));
  AOI21_X1  g605(.A(G176gat), .B1(new_n798_), .B2(new_n446_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(G1349gat));
  AOI21_X1  g607(.A(G183gat), .B1(new_n803_), .B2(new_n756_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n791_), .A2(new_n218_), .A3(new_n524_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1350gat));
  OAI21_X1  g610(.A(G190gat), .B1(new_n791_), .B2(new_n580_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n506_), .A2(new_n302_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n791_), .B2(new_n813_), .ZN(G1351gat));
  NAND3_X1  g613(.A1(new_n347_), .A2(new_n539_), .A3(new_n242_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT125), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n748_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n570_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(new_n480_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT126), .B(G197gat), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1352gat));
  NOR2_X1   g622(.A1(new_n820_), .A2(new_n445_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n247_), .A2(KEYINPUT127), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n247_), .A2(KEYINPUT127), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n824_), .B2(new_n825_), .ZN(G1353gat));
  AND2_X1   g627(.A1(new_n818_), .A2(new_n819_), .ZN(new_n829_));
  AOI211_X1 g628(.A(KEYINPUT63), .B(G211gat), .C1(new_n829_), .C2(new_n756_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT63), .B(G211gat), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n820_), .A2(new_n524_), .A3(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1354gat));
  AOI21_X1  g632(.A(G218gat), .B1(new_n829_), .B2(new_n506_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n829_), .A2(G218gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n510_), .B2(new_n835_), .ZN(G1355gat));
endmodule


