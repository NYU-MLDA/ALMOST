//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT85), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT84), .A2(KEYINPUT21), .ZN(new_n207_));
  AND2_X1   g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n206_), .B(new_n207_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G197gat), .A2(G204gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G197gat), .A2(G204gat), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n211_), .A2(KEYINPUT83), .A3(KEYINPUT21), .A4(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n208_), .A2(new_n209_), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT83), .B1(new_n216_), .B2(KEYINPUT21), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n203_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G218gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G211gat), .ZN(new_n220_));
  INV_X1    g019(.A(G211gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G218gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n211_), .A2(new_n212_), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT84), .A2(KEYINPUT21), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT84), .A2(KEYINPUT21), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n223_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n211_), .A2(KEYINPUT21), .A3(new_n212_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT83), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n228_), .A2(KEYINPUT85), .A3(new_n231_), .A4(new_n213_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n218_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT86), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(new_n229_), .B2(new_n214_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n223_), .A2(new_n216_), .A3(KEYINPUT86), .A4(KEYINPUT21), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G228gat), .ZN(new_n239_));
  INV_X1    g038(.A(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT29), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G155gat), .A2(G162gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT3), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G141gat), .A2(G148gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT2), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n245_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G141gat), .B(G148gat), .Z(new_n251_));
  NAND3_X1  g050(.A1(new_n244_), .A2(KEYINPUT81), .A3(KEYINPUT1), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(G155gat), .A3(G162gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n243_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT81), .B1(new_n244_), .B2(KEYINPUT1), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n251_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT82), .B(new_n251_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n250_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  OAI221_X1 g060(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .C1(new_n241_), .C2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT87), .B1(new_n261_), .B2(new_n241_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n250_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n260_), .ZN(new_n265_));
  AND2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n242_), .B1(new_n266_), .B2(new_n253_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n244_), .A2(KEYINPUT1), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT81), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(new_n270_), .A3(new_n252_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT82), .B1(new_n271_), .B2(new_n251_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n264_), .B1(new_n265_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT87), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT29), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n263_), .A2(new_n275_), .A3(new_n238_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n239_), .A2(new_n240_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n276_), .A2(KEYINPUT88), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT88), .B1(new_n276_), .B2(new_n277_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n262_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G78gat), .B(G106gat), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n261_), .A2(new_n241_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT28), .ZN(new_n284_));
  XOR2_X1   g083(.A(G22gat), .B(G50gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n281_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n287_), .B(new_n262_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n282_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n286_), .B1(new_n282_), .B2(new_n288_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT19), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT20), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n218_), .A2(new_n232_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT76), .ZN(new_n297_));
  INV_X1    g096(.A(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT23), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT25), .B(G183gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT26), .B(G190gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n304_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n302_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(KEYINPUT24), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n298_), .A2(KEYINPUT22), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT22), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G169gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n316_), .A3(new_n299_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n312_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n319_));
  INV_X1    g118(.A(G183gat), .ZN(new_n320_));
  INV_X1    g119(.A(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n318_), .A2(new_n319_), .B1(new_n306_), .B2(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n317_), .A2(new_n312_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT77), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n310_), .A2(new_n313_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n295_), .B1(new_n296_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT91), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n306_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n328_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n302_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(KEYINPUT91), .A3(new_n306_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n321_), .A2(KEYINPUT26), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n321_), .A2(KEYINPUT26), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT89), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT89), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n308_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n340_), .A3(new_n307_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n311_), .A2(new_n312_), .A3(new_n329_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n332_), .A2(new_n335_), .A3(new_n341_), .A4(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n306_), .A2(new_n322_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n324_), .A2(new_n344_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n343_), .A2(new_n345_), .B1(new_n233_), .B2(new_n237_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT92), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n327_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n335_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT91), .B1(new_n334_), .B2(new_n306_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n345_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n238_), .A3(new_n347_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n294_), .B1(new_n348_), .B2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n343_), .A2(new_n233_), .A3(new_n237_), .A4(new_n345_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n355_), .A2(KEYINPUT20), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT93), .ZN(new_n357_));
  INV_X1    g156(.A(new_n294_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n323_), .A2(new_n325_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n313_), .A2(new_n304_), .A3(new_n306_), .A4(new_n309_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n238_), .A2(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .A4(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n355_), .A3(KEYINPUT20), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT93), .B1(new_n364_), .B2(new_n294_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n354_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G8gat), .B(G36gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT18), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G64gat), .B(G92gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n354_), .A2(new_n363_), .A3(new_n365_), .A4(new_n370_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n373_), .A2(KEYINPUT27), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n351_), .A2(new_n238_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT92), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n379_), .A2(new_n358_), .A3(new_n352_), .A4(new_n327_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT98), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n347_), .B1(new_n351_), .B2(new_n238_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT20), .B1(new_n238_), .B2(new_n361_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n385_), .A2(KEYINPUT98), .A3(new_n358_), .A4(new_n352_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n364_), .A2(KEYINPUT97), .A3(new_n294_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT97), .B1(new_n364_), .B2(new_n294_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n371_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n377_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G1gat), .B(G29gat), .Z(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n395_), .B(new_n396_), .Z(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G127gat), .B(G134gat), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n399_), .A2(KEYINPUT79), .ZN(new_n400_));
  INV_X1    g199(.A(G134gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G127gat), .ZN(new_n402_));
  INV_X1    g201(.A(G127gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(G134gat), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n402_), .A2(new_n404_), .A3(KEYINPUT79), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G113gat), .B(G120gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n400_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n399_), .A2(KEYINPUT79), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n407_), .B1(new_n410_), .B2(new_n405_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n409_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(KEYINPUT80), .B(new_n407_), .C1(new_n410_), .C2(new_n405_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n273_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n409_), .A2(new_n411_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n261_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(KEYINPUT4), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n415_), .A2(new_n273_), .A3(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n419_), .A2(KEYINPUT94), .A3(new_n421_), .A4(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n416_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n421_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT94), .B1(new_n428_), .B2(new_n419_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n398_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT94), .ZN(new_n431_));
  INV_X1    g230(.A(new_n419_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(new_n427_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n433_), .A2(new_n397_), .A3(new_n425_), .A4(new_n424_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n376_), .A2(new_n392_), .A3(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n202_), .B1(new_n292_), .B2(new_n437_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n375_), .A2(new_n374_), .B1(new_n377_), .B2(new_n391_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n286_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n276_), .A2(new_n277_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n276_), .A2(KEYINPUT88), .A3(new_n277_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n287_), .B1(new_n445_), .B2(new_n262_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n288_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n440_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n289_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n439_), .A2(new_n449_), .A3(KEYINPUT99), .A4(new_n436_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n387_), .A2(new_n390_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n370_), .A2(KEYINPUT32), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(KEYINPUT96), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n354_), .A2(new_n363_), .A3(new_n365_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n435_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n434_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n426_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n459_), .A2(KEYINPUT33), .A3(new_n397_), .A4(new_n433_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n419_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n416_), .A2(new_n418_), .A3(new_n421_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n398_), .A3(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n372_), .A2(new_n373_), .A3(new_n464_), .ZN(new_n465_));
  OAI22_X1  g264(.A1(new_n453_), .A2(new_n456_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n292_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n438_), .A2(new_n450_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G227gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(G15gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n326_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT31), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G71gat), .B(G99gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G43gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n415_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n472_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n468_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n292_), .A2(new_n439_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n436_), .A2(new_n478_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT10), .B(G99gat), .Z(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G85gat), .B(G92gat), .Z(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT9), .ZN(new_n494_));
  INV_X1    g293(.A(G85gat), .ZN(new_n495_));
  INV_X1    g294(.A(G92gat), .ZN(new_n496_));
  OR3_X1    g295(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT9), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n489_), .A2(new_n492_), .A3(new_n494_), .A4(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  OR3_X1    g298(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n499_), .B(new_n500_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT8), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n501_), .A2(new_n493_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n501_), .B2(new_n493_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n498_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n508_));
  XOR2_X1   g307(.A(G71gat), .B(G78gat), .Z(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n508_), .A2(new_n509_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT12), .B1(new_n506_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n506_), .A2(new_n513_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n506_), .A2(KEYINPUT65), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT65), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n518_), .B(new_n498_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n517_), .A2(KEYINPUT12), .A3(new_n513_), .A4(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT66), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n516_), .A2(new_n520_), .A3(KEYINPUT66), .A4(new_n521_), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n506_), .B(new_n513_), .Z(new_n526_));
  OAI211_X1 g325(.A(new_n524_), .B(new_n525_), .C1(new_n521_), .C2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G120gat), .B(G148gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G176gat), .B(G204gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(new_n532_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n533_), .A2(KEYINPUT13), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT13), .B1(new_n533_), .B2(new_n534_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(G29gat), .B(G36gat), .Z(new_n539_));
  XOR2_X1   g338(.A(G43gat), .B(G50gat), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G29gat), .B(G36gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT73), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G1gat), .A2(G8gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT14), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G1gat), .B(G8gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT74), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n547_), .A2(new_n553_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n545_), .B(KEYINPUT15), .ZN(new_n561_));
  INV_X1    g360(.A(new_n553_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n563_), .A3(new_n558_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G169gat), .B(G197gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT75), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n565_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n538_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n485_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n545_), .B(new_n498_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT68), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT35), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n575_), .A2(KEYINPUT68), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n574_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n576_), .A2(KEYINPUT69), .A3(new_n583_), .A4(new_n581_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n517_), .A2(new_n561_), .A3(new_n519_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n579_), .A2(new_n580_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n582_), .A2(new_n584_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n589_), .B(KEYINPUT71), .Z(new_n591_));
  AND2_X1   g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n588_), .A2(new_n589_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT70), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(G134gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(G162gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n594_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n594_), .A2(new_n595_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n599_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n593_), .B2(KEYINPUT36), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT37), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n606_), .B(new_n600_), .C1(new_n601_), .C2(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n553_), .B(new_n609_), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(new_n513_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT72), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT17), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n613_), .B(new_n618_), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n611_), .A2(KEYINPUT17), .A3(new_n617_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n608_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n573_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT100), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n625_), .B1(new_n573_), .B2(new_n622_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n436_), .A2(G1gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT101), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n627_), .A2(new_n631_), .A3(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n537_), .A2(new_n621_), .A3(new_n570_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT102), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n485_), .A3(new_n604_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT103), .Z(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n435_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G1gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n630_), .A2(KEYINPUT38), .A3(new_n632_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n641_), .A3(new_n642_), .ZN(G1324gat));
  OAI21_X1  g442(.A(G8gat), .B1(new_n638_), .B2(new_n439_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT39), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n439_), .A2(G8gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n627_), .B2(new_n647_), .ZN(new_n648_));
  AND4_X1   g447(.A1(new_n646_), .A2(new_n624_), .A3(new_n626_), .A4(new_n647_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n645_), .B(KEYINPUT40), .C1(new_n648_), .C2(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  INV_X1    g453(.A(G15gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n639_), .B2(new_n478_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT41), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n623_), .A2(new_n655_), .A3(new_n478_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n639_), .B2(new_n449_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n623_), .A2(new_n660_), .A3(new_n449_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1327gat));
  INV_X1    g464(.A(new_n608_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n439_), .A2(new_n449_), .A3(new_n436_), .ZN(new_n667_));
  AOI22_X1  g466(.A1(new_n667_), .A2(new_n202_), .B1(new_n292_), .B2(new_n466_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n478_), .B1(new_n668_), .B2(new_n450_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n666_), .B1(new_n669_), .B2(new_n483_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n621_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT43), .B(new_n666_), .C1(new_n669_), .C2(new_n483_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n572_), .A4(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n483_), .B1(new_n468_), .B2(new_n479_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n675_), .B2(new_n608_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n621_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n676_), .A2(new_n673_), .A3(new_n677_), .A4(new_n572_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n674_), .A2(new_n680_), .A3(G29gat), .A4(new_n435_), .ZN(new_n681_));
  INV_X1    g480(.A(G29gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n604_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n677_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n572_), .B(new_n685_), .C1(new_n669_), .C2(new_n483_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n485_), .A2(KEYINPUT105), .A3(new_n572_), .A4(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n682_), .B1(new_n690_), .B2(new_n436_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n681_), .A2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(new_n439_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n674_), .A2(new_n680_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n439_), .A2(G36gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n688_), .A2(new_n689_), .A3(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT45), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT46), .Z(G1329gat));
  XNOR2_X1  g499(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n688_), .A2(new_n478_), .A3(new_n689_), .ZN(new_n704_));
  INV_X1    g503(.A(G43gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT106), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n708_), .A3(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n479_), .A2(new_n705_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n674_), .A2(new_n680_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n703_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n704_), .A2(new_n708_), .A3(new_n705_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n708_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n703_), .B(new_n712_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n702_), .B1(new_n713_), .B2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n712_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT108), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n716_), .A3(new_n701_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1330gat));
  NAND3_X1  g521(.A1(new_n674_), .A2(new_n680_), .A3(new_n449_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G50gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n292_), .A2(G50gat), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT109), .Z(new_n726_));
  OAI21_X1  g525(.A(new_n724_), .B1(new_n690_), .B2(new_n726_), .ZN(G1331gat));
  NOR2_X1   g526(.A1(new_n537_), .A2(new_n570_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n485_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n622_), .ZN(new_n730_));
  INV_X1    g529(.A(G57gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n435_), .ZN(new_n732_));
  AND4_X1   g531(.A1(new_n621_), .A2(new_n485_), .A3(new_n604_), .A4(new_n728_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(new_n435_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n734_), .B2(new_n731_), .ZN(G1332gat));
  INV_X1    g534(.A(G64gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n733_), .B2(new_n693_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT48), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n730_), .A2(new_n736_), .A3(new_n693_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n733_), .B2(new_n478_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n730_), .A2(new_n741_), .A3(new_n478_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1334gat));
  INV_X1    g545(.A(G78gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n733_), .B2(new_n449_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT50), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n730_), .A2(new_n747_), .A3(new_n449_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1335gat));
  NAND4_X1  g550(.A1(new_n676_), .A2(new_n673_), .A3(new_n677_), .A4(new_n728_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n436_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n729_), .A2(new_n684_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n495_), .A3(new_n435_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1336gat));
  OAI21_X1  g555(.A(G92gat), .B1(new_n752_), .B2(new_n439_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n754_), .A2(new_n496_), .A3(new_n693_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n752_), .B2(new_n479_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n754_), .A2(new_n490_), .A3(new_n478_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g562(.A(G106gat), .B1(new_n752_), .B2(new_n292_), .ZN(new_n764_));
  XOR2_X1   g563(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n765_));
  XNOR2_X1  g564(.A(new_n764_), .B(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n754_), .A2(new_n491_), .A3(new_n449_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1339gat));
  NOR3_X1   g570(.A1(new_n481_), .A2(new_n436_), .A3(new_n479_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n524_), .A2(new_n774_), .A3(new_n525_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n516_), .A2(new_n520_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(G230gat), .A3(G233gat), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n516_), .A2(new_n520_), .A3(KEYINPUT55), .A4(new_n521_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n773_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n779_), .B(KEYINPUT113), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n783_), .A2(KEYINPUT114), .A3(new_n775_), .A4(new_n777_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n785_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n532_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n570_), .A2(new_n533_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n785_), .B2(new_n532_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  INV_X1    g589(.A(new_n532_), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n790_), .B(new_n791_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n789_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n788_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n568_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n565_), .A2(new_n796_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n554_), .A2(new_n563_), .A3(new_n559_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n557_), .A2(new_n558_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n796_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n800_), .B2(KEYINPUT116), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n802_), .A3(new_n796_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n797_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n533_), .A2(new_n534_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n604_), .B1(new_n795_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n804_), .A2(new_n533_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n608_), .B1(new_n811_), .B2(new_n810_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n807_), .A2(new_n808_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT57), .B(new_n604_), .C1(new_n795_), .C2(new_n806_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n621_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n608_), .A2(new_n621_), .A3(new_n571_), .A4(new_n537_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n817_), .B(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT59), .B(new_n772_), .C1(new_n816_), .C2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n785_), .A2(new_n532_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n790_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n532_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n794_), .A3(new_n824_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n786_), .A2(new_n787_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n806_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n808_), .B1(new_n827_), .B2(new_n683_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n813_), .A2(new_n812_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n815_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n819_), .B1(new_n830_), .B2(new_n677_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n772_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n821_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n820_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n571_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n830_), .A2(new_n677_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n819_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n772_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n571_), .A2(G113gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n836_), .B1(new_n840_), .B2(new_n841_), .ZN(G1340gat));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n834_), .B2(new_n538_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n537_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(KEYINPUT60), .B2(new_n843_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n840_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT117), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n537_), .B1(new_n820_), .B2(new_n833_), .ZN(new_n850_));
  OAI221_X1 g649(.A(new_n849_), .B1(new_n840_), .B2(new_n846_), .C1(new_n850_), .C2(new_n843_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(G1341gat));
  OAI21_X1  g651(.A(G127gat), .B1(new_n835_), .B2(new_n677_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n621_), .A2(new_n403_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n840_), .B2(new_n854_), .ZN(G1342gat));
  OAI21_X1  g654(.A(G134gat), .B1(new_n835_), .B2(new_n608_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n683_), .A2(new_n401_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n840_), .B2(new_n857_), .ZN(G1343gat));
  NOR4_X1   g657(.A1(new_n693_), .A2(new_n292_), .A3(new_n436_), .A4(new_n478_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n839_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n570_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n538_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g664(.A1(new_n860_), .A2(new_n677_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT61), .B(G155gat), .Z(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  OR3_X1    g667(.A1(new_n860_), .A2(G162gat), .A3(new_n604_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G162gat), .B1(new_n860_), .B2(new_n608_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1347gat));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n439_), .A2(new_n449_), .A3(new_n482_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n839_), .A2(new_n570_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n874_), .B2(G169gat), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n839_), .A2(new_n873_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n570_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT119), .Z(new_n879_));
  AOI22_X1  g678(.A1(new_n875_), .A2(new_n876_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n875_), .A2(new_n876_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n874_), .A2(new_n872_), .A3(G169gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(G1348gat));
  NAND2_X1  g682(.A1(new_n877_), .A2(new_n538_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g684(.A1(new_n877_), .A2(new_n621_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT120), .B1(new_n886_), .B2(new_n307_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n320_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889_));
  INV_X1    g688(.A(new_n307_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n877_), .A2(new_n889_), .A3(new_n621_), .A4(new_n890_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n887_), .A2(new_n888_), .A3(new_n891_), .ZN(G1350gat));
  NAND4_X1  g691(.A1(new_n877_), .A2(new_n683_), .A3(new_n338_), .A4(new_n340_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n877_), .A2(new_n666_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n321_), .ZN(G1351gat));
  NAND3_X1  g694(.A1(new_n449_), .A2(new_n436_), .A3(new_n479_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n896_), .A2(KEYINPUT121), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(KEYINPUT121), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n897_), .A2(new_n693_), .A3(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n831_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n570_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT122), .B(G197gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1352gat));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n538_), .ZN(new_n905_));
  INV_X1    g704(.A(G204gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(KEYINPUT123), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n905_), .B(new_n907_), .ZN(G1353gat));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n621_), .B1(new_n909_), .B2(new_n221_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT124), .Z(new_n911_));
  NAND2_X1  g710(.A1(new_n901_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n221_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1354gat));
  XOR2_X1   g713(.A(KEYINPUT126), .B(G218gat), .Z(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n683_), .B(new_n899_), .C1(new_n816_), .C2(new_n819_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n901_), .A2(KEYINPUT125), .A3(new_n683_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n916_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n901_), .A2(new_n666_), .A3(new_n916_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(KEYINPUT127), .B1(new_n921_), .B2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(KEYINPUT125), .B1(new_n901_), .B2(new_n683_), .ZN(new_n925_));
  NOR4_X1   g724(.A1(new_n831_), .A2(new_n918_), .A3(new_n604_), .A4(new_n900_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n915_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(new_n928_), .A3(new_n922_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n924_), .A2(new_n929_), .ZN(G1355gat));
endmodule


