//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G71gat), .B(G78gat), .ZN(new_n205_));
  OR3_X1    g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n202_), .A2(new_n205_), .A3(KEYINPUT11), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR3_X1   g010(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n209_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT6), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT67), .A3(new_n210_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n215_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G85gat), .B(G92gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT68), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(KEYINPUT68), .A3(new_n221_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT8), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT69), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n215_), .A2(new_n210_), .A3(new_n218_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n221_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n224_), .A2(KEYINPUT69), .A3(KEYINPUT8), .A4(new_n225_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n215_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n235_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n237_));
  INV_X1    g036(.A(G85gat), .ZN(new_n238_));
  INV_X1    g037(.A(G92gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT9), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT65), .ZN(new_n242_));
  OAI22_X1  g041(.A1(new_n240_), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n236_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n234_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT10), .B(G99gat), .ZN(new_n247_));
  OAI221_X1 g046(.A(new_n246_), .B1(new_n245_), .B2(new_n244_), .C1(G106gat), .C2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n208_), .B1(new_n233_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT12), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n233_), .A2(new_n248_), .A3(new_n208_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G230gat), .A2(G233gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n253_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n251_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n233_), .A2(KEYINPUT70), .A3(new_n248_), .A4(new_n208_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n233_), .A2(new_n248_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n208_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n254_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n257_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G120gat), .B(G148gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(G204gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT5), .B(G176gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n270_), .B(new_n271_), .Z(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n272_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n257_), .A2(new_n267_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT13), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n273_), .A2(KEYINPUT13), .A3(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n278_), .A2(KEYINPUT72), .A3(new_n279_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G15gat), .B(G22gat), .ZN(new_n285_));
  INV_X1    g084(.A(G1gat), .ZN(new_n286_));
  INV_X1    g085(.A(G8gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT14), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G1gat), .B(G8gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G29gat), .B(G36gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(G43gat), .B(G50gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n291_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT78), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G229gat), .A2(G233gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n294_), .B(KEYINPUT15), .Z(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n291_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n294_), .B2(new_n291_), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n297_), .B(KEYINPUT79), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G113gat), .B(G141gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G169gat), .B(G197gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n305_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n284_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n208_), .B(new_n291_), .Z(new_n312_));
  NAND2_X1  g111(.A1(G231gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G183gat), .B(G211gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G127gat), .B(G155gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT17), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n319_), .B(KEYINPUT17), .Z(new_n322_));
  OAI21_X1  g121(.A(new_n321_), .B1(new_n314_), .B2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT77), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G8gat), .B(G36gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(G92gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT18), .B(G64gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  NOR2_X1   g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT24), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G183gat), .ZN(new_n335_));
  OR3_X1    g134(.A1(new_n335_), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT26), .B(G190gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT25), .B1(new_n335_), .B2(KEYINPUT80), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n332_), .A2(KEYINPUT24), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n334_), .A2(KEYINPUT82), .A3(new_n339_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT23), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .A4(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(G183gat), .B2(G190gat), .ZN(new_n348_));
  INV_X1    g147(.A(G169gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT22), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT83), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n353_));
  INV_X1    g152(.A(G176gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT22), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G169gat), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .A4(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n348_), .A2(new_n333_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n347_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G197gat), .B(G204gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT21), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G211gat), .B(G218gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n362_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n363_), .A2(new_n364_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n360_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n369_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n330_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n346_), .B1(KEYINPUT24), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT92), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT25), .B(G183gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n337_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(new_n377_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n378_), .A2(new_n334_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n356_), .A2(new_n350_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n333_), .B1(new_n383_), .B2(G176gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT93), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n348_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n374_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n371_), .A2(KEYINPUT20), .A3(new_n373_), .A4(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT20), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n359_), .B2(new_n374_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n374_), .A2(new_n387_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n373_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n329_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G141gat), .A2(G148gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G141gat), .ZN(new_n399_));
  INV_X1    g198(.A(G148gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n398_), .B1(KEYINPUT3), .B2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n401_), .A2(KEYINPUT3), .ZN(new_n403_));
  NOR2_X1   g202(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT87), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G155gat), .B(G162gat), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n408_), .A2(KEYINPUT88), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT87), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n402_), .A2(new_n403_), .A3(new_n410_), .A4(new_n405_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(KEYINPUT88), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n407_), .A2(new_n409_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(G155gat), .A2(G162gat), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n414_), .A2(KEYINPUT1), .B1(new_n399_), .B2(new_n400_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n415_), .B(new_n396_), .C1(KEYINPUT1), .C2(new_n408_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G127gat), .B(G134gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G113gat), .B(G120gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n418_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT94), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT95), .Z(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n413_), .A2(new_n416_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n421_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n417_), .A2(new_n422_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n423_), .B(new_n427_), .C1(new_n431_), .C2(new_n418_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n431_), .A2(new_n425_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(new_n238_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT0), .B(G57gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n432_), .A2(new_n433_), .A3(KEYINPUT33), .A4(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n329_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n392_), .A2(new_n393_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n389_), .B(new_n440_), .C1(new_n441_), .C2(new_n373_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n395_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n423_), .B1(new_n431_), .B2(new_n418_), .ZN(new_n444_));
  OAI22_X1  g243(.A1(new_n444_), .A2(new_n425_), .B1(new_n431_), .B2(new_n426_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n438_), .B1(new_n445_), .B2(KEYINPUT33), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n432_), .A2(new_n433_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n437_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n432_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n389_), .B1(new_n441_), .B2(new_n373_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n329_), .A2(KEYINPUT32), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n451_), .A2(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n371_), .A2(KEYINPUT20), .A3(new_n388_), .ZN(new_n456_));
  MUX2_X1   g255(.A(new_n456_), .B(new_n441_), .S(new_n373_), .Z(new_n457_));
  OR2_X1    g256(.A1(new_n457_), .A2(new_n454_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n447_), .A2(new_n450_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n359_), .A2(KEYINPUT30), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT30), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n347_), .B2(new_n358_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT85), .B1(new_n460_), .B2(new_n462_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT31), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT84), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G15gat), .B(G43gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G71gat), .B(G99gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n466_), .A2(new_n467_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n467_), .B1(new_n466_), .B2(new_n474_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n476_), .A2(new_n421_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n360_), .A2(new_n461_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n462_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n464_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT31), .B1(new_n481_), .B2(new_n473_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n422_), .B1(new_n482_), .B2(new_n475_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n465_), .B1(new_n478_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n421_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n465_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n422_), .A3(new_n475_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G228gat), .A2(G233gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n492_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n370_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n417_), .A2(KEYINPUT29), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(new_n490_), .A3(new_n374_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G78gat), .B(G106gat), .Z(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n497_), .B(new_n499_), .ZN(new_n500_));
  OR3_X1    g299(.A1(new_n417_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(G50gat), .B1(new_n417_), .B2(KEYINPUT29), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT28), .B(G22gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(new_n504_), .A3(new_n502_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n500_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n497_), .A2(KEYINPUT90), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n494_), .A2(new_n496_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n498_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  OAI22_X1  g312(.A1(new_n513_), .A2(KEYINPUT91), .B1(new_n497_), .B2(new_n499_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n506_), .A2(new_n507_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n494_), .A2(new_n496_), .A3(new_n511_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n511_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n499_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n515_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n509_), .B1(new_n514_), .B2(new_n520_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n459_), .A2(new_n489_), .A3(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(KEYINPUT27), .B(new_n395_), .C1(new_n457_), .C2(new_n329_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n395_), .A2(new_n442_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(KEYINPUT27), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n508_), .B1(new_n513_), .B2(KEYINPUT91), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n497_), .A2(new_n499_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n526_), .A2(new_n528_), .B1(new_n500_), .B2(new_n508_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n488_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n486_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n521_), .A2(new_n488_), .A3(new_n484_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n525_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n451_), .A2(new_n452_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n522_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n311_), .A2(new_n325_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT74), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT34), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n262_), .A2(new_n299_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n546_), .B(new_n547_), .C1(new_n294_), .C2(new_n262_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n545_), .A2(new_n541_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n549_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(G162gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT73), .B(G134gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT36), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n550_), .A2(new_n551_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n555_), .A2(KEYINPUT36), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n540_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(new_n539_), .A3(new_n558_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n538_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n286_), .A3(new_n535_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT38), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n571_), .A2(KEYINPUT96), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n569_), .A2(new_n570_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(KEYINPUT96), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n563_), .A2(new_n558_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n538_), .A2(new_n535_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(G1gat), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .A4(new_n578_), .ZN(G1324gat));
  NAND3_X1  g378(.A1(new_n538_), .A2(new_n576_), .A3(new_n525_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT97), .B(KEYINPUT39), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n580_), .A2(G8gat), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n580_), .B2(G8gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n525_), .A2(new_n287_), .ZN(new_n584_));
  OAI22_X1  g383(.A1(new_n582_), .A2(new_n583_), .B1(new_n567_), .B2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g385(.A(new_n489_), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n567_), .A2(G15gat), .A3(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n538_), .A2(new_n576_), .A3(new_n489_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(G15gat), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT98), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT41), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(KEYINPUT98), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n592_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n588_), .B1(new_n594_), .B2(new_n595_), .ZN(G1326gat));
  OR3_X1    g395(.A1(new_n567_), .A2(G22gat), .A3(new_n529_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n538_), .A2(new_n576_), .A3(new_n521_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT99), .B(KEYINPUT42), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n598_), .A2(G22gat), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n598_), .B2(G22gat), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(G1327gat));
  INV_X1    g401(.A(new_n537_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n575_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n282_), .A2(new_n283_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n606_), .A2(new_n309_), .A3(new_n324_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(G29gat), .B1(new_n609_), .B2(new_n535_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT43), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n565_), .B2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n537_), .B2(new_n566_), .ZN(new_n614_));
  AOI211_X1 g413(.A(new_n535_), .B(new_n525_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n615_));
  OAI221_X1 g414(.A(new_n565_), .B1(new_n612_), .B2(new_n611_), .C1(new_n615_), .C2(new_n522_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n607_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT44), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT101), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n621_));
  AOI211_X1 g420(.A(new_n621_), .B(KEYINPUT44), .C1(new_n617_), .C2(new_n607_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n617_), .A2(KEYINPUT44), .A3(new_n607_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n625_), .A2(G29gat), .A3(new_n535_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n610_), .B1(new_n624_), .B2(new_n626_), .ZN(G1328gat));
  INV_X1    g426(.A(new_n525_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n608_), .A2(G36gat), .A3(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT45), .Z(new_n630_));
  OAI211_X1 g429(.A(new_n525_), .B(new_n625_), .C1(new_n620_), .C2(new_n622_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n631_), .A2(new_n632_), .A3(G36gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n631_), .B2(G36gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT46), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT46), .B(new_n630_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1329gat));
  AOI21_X1  g438(.A(G43gat), .B1(new_n609_), .B2(new_n489_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n489_), .A2(G43gat), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n623_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n640_), .B1(new_n642_), .B2(new_n625_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g443(.A1(new_n625_), .A2(G50gat), .A3(new_n521_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n608_), .A2(new_n529_), .ZN(new_n646_));
  OAI22_X1  g445(.A1(new_n645_), .A2(new_n623_), .B1(G50gat), .B2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT103), .Z(G1331gat));
  NOR2_X1   g447(.A1(new_n284_), .A2(new_n325_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n566_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT104), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n537_), .A2(new_n310_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(KEYINPUT104), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(G57gat), .A3(new_n536_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n649_), .A2(new_n576_), .A3(new_n652_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT105), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n535_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n655_), .B1(new_n658_), .B2(G57gat), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1332gat));
  OR3_X1    g460(.A1(new_n654_), .A2(G64gat), .A3(new_n628_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n657_), .A2(new_n525_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n663_), .A2(G64gat), .A3(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n663_), .B2(G64gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n665_), .B2(new_n666_), .ZN(G1333gat));
  NAND2_X1  g466(.A1(new_n657_), .A2(new_n489_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT49), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(new_n669_), .A3(G71gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n668_), .B2(G71gat), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n587_), .A2(G71gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT108), .ZN(new_n673_));
  OAI22_X1  g472(.A1(new_n670_), .A2(new_n671_), .B1(new_n654_), .B2(new_n673_), .ZN(G1334gat));
  INV_X1    g473(.A(KEYINPUT50), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n657_), .A2(new_n521_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(G78gat), .ZN(new_n677_));
  INV_X1    g476(.A(G78gat), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT50), .B(new_n678_), .C1(new_n657_), .C2(new_n521_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n521_), .A2(new_n678_), .ZN(new_n680_));
  OAI22_X1  g479(.A1(new_n677_), .A2(new_n679_), .B1(new_n654_), .B2(new_n680_), .ZN(G1335gat));
  NOR3_X1   g480(.A1(new_n284_), .A2(new_n310_), .A3(new_n324_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n605_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n238_), .A3(new_n535_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n617_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT109), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT109), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n536_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n689_), .B2(new_n238_), .ZN(G1336gat));
  NAND3_X1  g489(.A1(new_n684_), .A2(new_n239_), .A3(new_n525_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n628_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(new_n239_), .ZN(G1337gat));
  NOR3_X1   g492(.A1(new_n683_), .A2(new_n247_), .A3(new_n587_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n682_), .A2(new_n617_), .A3(new_n489_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(G99gat), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT51), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT111), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n696_), .B(new_n699_), .ZN(G1338gat));
  NAND3_X1  g499(.A1(new_n682_), .A2(new_n617_), .A3(new_n521_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT112), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n702_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(G106gat), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT52), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT52), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n703_), .A2(new_n707_), .A3(G106gat), .A4(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  OR3_X1    g508(.A1(new_n683_), .A2(G106gat), .A3(new_n529_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT53), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT53), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n713_), .A3(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1339gat));
  NOR2_X1   g514(.A1(new_n525_), .A2(new_n536_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n532_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT115), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(KEYINPUT58), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n264_), .A2(new_n250_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n249_), .A2(KEYINPUT12), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n261_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n266_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT114), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT55), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n256_), .A2(new_n255_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n722_), .A2(new_n723_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n251_), .B(KEYINPUT55), .C1(new_n255_), .C2(new_n256_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT114), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n724_), .A2(new_n732_), .A3(new_n266_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n726_), .A2(new_n730_), .A3(new_n731_), .A4(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT56), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n272_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n734_), .B2(new_n272_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n275_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n298_), .A2(new_n304_), .A3(new_n308_), .ZN(new_n740_));
  MUX2_X1   g539(.A(new_n301_), .B(new_n296_), .S(new_n302_), .Z(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n308_), .B2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n721_), .B1(new_n739_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n734_), .A2(new_n272_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT56), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n734_), .A2(new_n735_), .A3(new_n272_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n745_), .A2(new_n275_), .A3(new_n742_), .A4(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n721_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n565_), .B1(new_n743_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT116), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n745_), .A2(new_n310_), .A3(new_n275_), .A4(new_n746_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n276_), .A2(new_n742_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT57), .B1(new_n755_), .B2(new_n576_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT57), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n757_), .B(new_n575_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT116), .B(new_n565_), .C1(new_n743_), .C2(new_n749_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n752_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n325_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n278_), .A2(new_n309_), .A3(new_n279_), .A4(new_n324_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n765_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n763_), .B1(new_n768_), .B2(new_n566_), .ZN(new_n769_));
  AOI211_X1 g568(.A(KEYINPUT54), .B(new_n565_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n719_), .B1(new_n762_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT117), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n771_), .B1(new_n761_), .B2(new_n325_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n719_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(G113gat), .B1(new_n778_), .B2(new_n310_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT59), .B1(new_n776_), .B2(new_n719_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n324_), .B1(new_n759_), .B2(new_n750_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n781_), .B(new_n718_), .C1(new_n782_), .C2(new_n771_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(G113gat), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(new_n309_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n779_), .A2(new_n786_), .ZN(G1340gat));
  OAI211_X1 g586(.A(new_n606_), .B(new_n783_), .C1(new_n773_), .C2(new_n781_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT119), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n780_), .A2(new_n790_), .A3(new_n606_), .A4(new_n783_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n789_), .A2(G120gat), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(G120gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n284_), .B2(KEYINPUT60), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT118), .B1(new_n793_), .B2(KEYINPUT60), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n778_), .B(new_n796_), .C1(new_n797_), .C2(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n792_), .A2(new_n798_), .ZN(G1341gat));
  NAND2_X1  g598(.A1(new_n778_), .A2(new_n324_), .ZN(new_n800_));
  INV_X1    g599(.A(G127gat), .ZN(new_n801_));
  NOR2_X1   g600(.A1(KEYINPUT120), .A2(G127gat), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n784_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(G127gat), .B1(new_n325_), .B2(KEYINPUT120), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n800_), .A2(new_n801_), .B1(new_n803_), .B2(new_n804_), .ZN(G1342gat));
  AOI21_X1  g604(.A(G134gat), .B1(new_n778_), .B2(new_n575_), .ZN(new_n806_));
  INV_X1    g605(.A(G134gat), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n784_), .A2(new_n807_), .A3(new_n566_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1343gat));
  NOR2_X1   g608(.A1(new_n776_), .A2(new_n533_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n310_), .A3(new_n716_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(KEYINPUT121), .B(G141gat), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n811_), .B(new_n812_), .Z(G1344gat));
  NAND3_X1  g612(.A1(new_n810_), .A2(new_n606_), .A3(new_n716_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g614(.A1(new_n810_), .A2(new_n324_), .A3(new_n716_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT61), .B(G155gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1346gat));
  AND2_X1   g617(.A1(new_n565_), .A2(G162gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n810_), .A2(new_n716_), .A3(new_n819_), .ZN(new_n820_));
  NOR4_X1   g619(.A1(new_n776_), .A2(new_n576_), .A3(new_n533_), .A4(new_n717_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(G162gat), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT122), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n820_), .B(new_n824_), .C1(G162gat), .C2(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1347gat));
  NOR2_X1   g625(.A1(new_n628_), .A2(new_n535_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n532_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n310_), .B(new_n829_), .C1(new_n782_), .C2(new_n771_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G169gat), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n831_), .A2(KEYINPUT124), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(KEYINPUT124), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n833_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n831_), .A2(KEYINPUT124), .A3(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n835_), .B(new_n837_), .C1(new_n383_), .C2(new_n830_), .ZN(G1348gat));
  OAI21_X1  g637(.A(new_n829_), .B1(new_n782_), .B2(new_n771_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G176gat), .B1(new_n840_), .B2(new_n606_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n829_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n776_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n284_), .A2(new_n354_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(G1349gat));
  OR3_X1    g644(.A1(new_n839_), .A2(new_n325_), .A3(new_n379_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n776_), .A2(new_n325_), .A3(new_n842_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(G183gat), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT125), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n846_), .B(KEYINPUT125), .C1(G183gat), .C2(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1350gat));
  OAI21_X1  g651(.A(G190gat), .B1(new_n839_), .B2(new_n566_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n575_), .A2(new_n337_), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT126), .Z(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n839_), .B2(new_n855_), .ZN(G1351gat));
  NOR3_X1   g655(.A1(new_n776_), .A2(new_n533_), .A3(new_n828_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n310_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n606_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n324_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT63), .B(G211gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n862_), .B2(new_n865_), .ZN(G1354gat));
  AOI21_X1  g665(.A(G218gat), .B1(new_n857_), .B2(new_n575_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n565_), .A2(G218gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n857_), .B2(new_n868_), .ZN(G1355gat));
endmodule


