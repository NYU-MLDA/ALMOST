//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(KEYINPUT82), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT82), .ZN(new_n205_));
  NAND4_X1  g004(.A1(new_n205_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(KEYINPUT82), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .A4(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT83), .B1(new_n209_), .B2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n206_), .A2(new_n208_), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n205_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n205_), .A2(KEYINPUT2), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT83), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .A4(new_n212_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT81), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n214_), .A2(new_n220_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n202_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n224_), .B(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n229_), .B1(G141gat), .B2(G148gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n225_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(KEYINPUT4), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G225gat), .A2(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n231_), .A2(new_n241_), .A3(new_n235_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n236_), .A2(KEYINPUT91), .A3(new_n239_), .A4(new_n237_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n236_), .A2(new_n239_), .A3(new_n237_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT91), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G1gat), .B(G29gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G85gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT0), .B(G57gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT97), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n248_), .A2(new_n252_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n248_), .A2(KEYINPUT97), .A3(new_n252_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G226gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT19), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n261_));
  OR2_X1    g060(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n263_));
  AOI21_X1  g062(.A(G176gat), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n261_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n263_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(KEYINPUT80), .A3(new_n265_), .ZN(new_n272_));
  INV_X1    g071(.A(G183gat), .ZN(new_n273_));
  INV_X1    g072(.A(G190gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT23), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(G183gat), .A3(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n274_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n267_), .A2(new_n272_), .A3(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G190gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n273_), .A2(KEYINPUT25), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT77), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT25), .B(G183gat), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n282_), .B(new_n285_), .C1(new_n286_), .C2(new_n284_), .ZN(new_n287_));
  INV_X1    g086(.A(G169gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n268_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(KEYINPUT24), .A3(new_n265_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(KEYINPUT78), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n277_), .A2(KEYINPUT79), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT79), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n293_), .A2(new_n276_), .A3(G183gat), .A4(G190gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n275_), .A3(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n289_), .A2(KEYINPUT24), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n287_), .A2(new_n290_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n281_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G197gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n305_));
  INV_X1    g104(.A(G204gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n305_), .B1(G197gat), .B2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(G197gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n304_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G211gat), .B(G218gat), .Z(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(KEYINPUT21), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT21), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n313_), .B(new_n304_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n310_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n303_), .A2(G204gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT21), .B1(new_n308_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT86), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n314_), .A2(new_n315_), .A3(KEYINPUT86), .A4(new_n317_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n312_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT20), .B1(new_n302_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n282_), .A2(new_n286_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n297_), .A2(new_n278_), .A3(new_n290_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n295_), .A2(new_n279_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n264_), .A2(new_n266_), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n324_), .A2(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT95), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI211_X1 g129(.A(new_n266_), .B(new_n264_), .C1(new_n295_), .C2(new_n279_), .ZN(new_n331_));
  AND4_X1   g130(.A1(new_n278_), .A2(new_n324_), .A3(new_n290_), .A4(new_n297_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT95), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n330_), .A2(new_n322_), .A3(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n260_), .B1(new_n323_), .B2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n260_), .B(KEYINPUT88), .Z(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n320_), .A2(new_n321_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n311_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n328_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n299_), .A2(new_n300_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n342_), .A2(new_n297_), .A3(new_n291_), .A4(new_n295_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n281_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n322_), .A3(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n345_), .A3(KEYINPUT20), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n335_), .B1(new_n337_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT96), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G64gat), .B(G92gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  AND2_X1   g152(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n347_), .A2(new_n348_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT20), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n356_), .B1(new_n302_), .B2(new_n322_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n336_), .B1(new_n357_), .B2(new_n341_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n260_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n323_), .A2(new_n360_), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n358_), .A2(new_n361_), .A3(new_n354_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n347_), .A2(new_n354_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT96), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n258_), .A2(new_n355_), .A3(new_n362_), .A4(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n353_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT90), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n346_), .A2(new_n337_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n290_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT77), .B1(new_n273_), .B2(KEYINPUT25), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(G183gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n283_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n374_), .B2(KEYINPUT77), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n370_), .B1(new_n375_), .B2(new_n282_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n297_), .B1(new_n376_), .B2(KEYINPUT78), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n291_), .A2(new_n295_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n344_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n356_), .B1(new_n379_), .B2(new_n339_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n260_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n369_), .A2(new_n353_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n367_), .A2(new_n368_), .A3(new_n383_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n346_), .A2(new_n337_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(KEYINPUT90), .A3(new_n353_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(KEYINPUT92), .B(KEYINPUT33), .Z(new_n388_));
  NAND2_X1  g187(.A1(new_n256_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n236_), .A2(new_n240_), .A3(new_n237_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n252_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT93), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n238_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT93), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n394_), .A3(new_n252_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT94), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n392_), .A2(KEYINPUT94), .A3(new_n393_), .A4(new_n395_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n248_), .A2(new_n252_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT92), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(KEYINPUT33), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n387_), .A2(new_n389_), .A3(new_n400_), .A4(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n365_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI211_X1 g208(.A(KEYINPUT30), .B(new_n281_), .C1(new_n296_), .C2(new_n301_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n235_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n379_), .A2(KEYINPUT30), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n343_), .A2(new_n411_), .A3(new_n344_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n234_), .A3(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G15gat), .B(G43gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT31), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n413_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n409_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n410_), .A2(new_n412_), .A3(new_n235_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n234_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n418_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n413_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n408_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G106gat), .ZN(new_n430_));
  AOI211_X1 g229(.A(new_n210_), .B(new_n226_), .C1(new_n223_), .C2(new_n228_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n215_), .A2(new_n218_), .A3(new_n212_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n432_), .A2(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n223_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n209_), .A2(new_n213_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n435_), .B2(new_n219_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n431_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n339_), .B(new_n430_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G228gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(G78gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n438_), .B1(new_n225_), .B2(new_n230_), .ZN(new_n443_));
  OAI21_X1  g242(.A(G106gat), .B1(new_n443_), .B2(new_n322_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n439_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n442_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT87), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n442_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n231_), .A2(KEYINPUT29), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n430_), .B1(new_n449_), .B2(new_n339_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n443_), .A2(new_n322_), .A3(G106gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n448_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n439_), .A2(new_n444_), .A3(new_n442_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n437_), .A2(new_n438_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G22gat), .B(G50gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n456_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n447_), .A2(new_n455_), .A3(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n460_), .B(KEYINPUT87), .C1(new_n445_), .C2(new_n446_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n429_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n428_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n462_), .A2(new_n422_), .A3(new_n427_), .A4(new_n463_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n258_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n330_), .A2(new_n333_), .A3(new_n322_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n359_), .B1(new_n380_), .B2(new_n470_), .ZN(new_n471_));
  AND4_X1   g270(.A1(KEYINPUT20), .A2(new_n341_), .A3(new_n345_), .A4(new_n336_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n366_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT98), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT98), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n347_), .A2(new_n475_), .A3(new_n366_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT27), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n385_), .B2(new_n353_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(KEYINPUT99), .B(KEYINPUT27), .Z(new_n480_));
  NAND3_X1  g279(.A1(new_n384_), .A2(new_n386_), .A3(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n405_), .A2(new_n466_), .B1(new_n469_), .B2(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G15gat), .B(G22gat), .Z(new_n484_));
  NAND2_X1  g283(.A1(G1gat), .A2(G8gat), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(KEYINPUT14), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT75), .ZN(new_n487_));
  XOR2_X1   g286(.A(G1gat), .B(G8gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT75), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n486_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n488_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G43gat), .B(G50gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(G29gat), .B(G36gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n498_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n494_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(KEYINPUT76), .A3(new_n501_), .ZN(new_n502_));
  OR3_X1    g301(.A1(new_n494_), .A2(KEYINPUT76), .A3(new_n500_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n502_), .A2(G229gat), .A3(G233gat), .A4(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n498_), .B(KEYINPUT15), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n495_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n501_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G169gat), .B(G197gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n504_), .A2(new_n508_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G57gat), .B(G64gat), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(KEYINPUT11), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(KEYINPUT11), .ZN(new_n520_));
  XOR2_X1   g319(.A(G71gat), .B(G78gat), .Z(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n520_), .A2(new_n521_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT67), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G85gat), .B(G92gat), .Z(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT10), .B(G99gat), .Z(new_n529_));
  AOI22_X1  g328(.A1(KEYINPUT9), .A2(new_n528_), .B1(new_n529_), .B2(new_n430_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(KEYINPUT9), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT6), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT64), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT64), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT6), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n534_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n530_), .A2(new_n532_), .A3(new_n536_), .A4(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT7), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n542_), .A3(new_n536_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n546_), .A2(new_n528_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n547_), .B1(new_n546_), .B2(new_n528_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n543_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT66), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(KEYINPUT66), .B(new_n543_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n527_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n551_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n553_), .A3(new_n526_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(G230gat), .A3(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n550_), .A2(KEYINPUT12), .A3(new_n523_), .A4(new_n522_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n561_), .A2(new_n555_), .A3(new_n562_), .A4(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G120gat), .B(G148gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(G204gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT5), .B(G176gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n559_), .A2(new_n564_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT13), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n569_), .B1(new_n559_), .B2(new_n564_), .ZN(new_n573_));
  OR3_X1    g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n483_), .A2(new_n517_), .A3(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n500_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT34), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT68), .B(KEYINPUT35), .Z(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n580_), .A2(new_n581_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n505_), .A2(new_n550_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n578_), .A2(new_n582_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n498_), .B1(new_n556_), .B2(new_n553_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n584_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n580_), .B(new_n581_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G134gat), .B(G162gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n585_), .A2(new_n587_), .A3(new_n590_), .A4(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT74), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n585_), .A2(new_n590_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n595_), .B(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n597_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n600_), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT74), .B(new_n602_), .C1(new_n585_), .C2(new_n590_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n596_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n602_), .B1(new_n585_), .B2(new_n590_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT73), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(KEYINPUT73), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n608_), .A2(KEYINPUT37), .A3(new_n596_), .A4(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n494_), .B(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n614_), .A2(new_n524_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n524_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(G211gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT16), .B(G183gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT17), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT67), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n617_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n615_), .A2(KEYINPUT67), .A3(new_n616_), .A4(new_n622_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n621_), .A2(KEYINPUT17), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n612_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n577_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n258_), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n630_), .A2(G1gat), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT102), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n632_), .A2(new_n633_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(KEYINPUT102), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n604_), .A2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT100), .B(new_n596_), .C1(new_n601_), .C2(new_n603_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT101), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n640_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n627_), .A3(new_n577_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n631_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .A4(new_n648_), .ZN(G1324gat));
  OAI21_X1  g448(.A(G8gat), .B1(new_n647_), .B2(new_n482_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT39), .ZN(new_n651_));
  OR3_X1    g450(.A1(new_n630_), .A2(G8gat), .A3(new_n482_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT40), .ZN(G1325gat));
  OR3_X1    g453(.A1(new_n630_), .A2(G15gat), .A3(new_n429_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n647_), .A2(new_n429_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(G15gat), .A3(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n656_), .B2(G15gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT104), .ZN(G1326gat));
  OR3_X1    g460(.A1(new_n630_), .A2(G22gat), .A3(new_n464_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G22gat), .B1(new_n647_), .B2(new_n464_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT105), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n666_), .B(G22gat), .C1(new_n647_), .C2(new_n464_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n664_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n665_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n662_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(G1327gat));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n467_), .A2(new_n468_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n674_), .A2(new_n631_), .A3(new_n482_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n465_), .B1(new_n365_), .B2(new_n404_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n673_), .B(new_n611_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT107), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n483_), .B2(new_n612_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n405_), .A2(new_n466_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n469_), .A2(new_n482_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n673_), .A4(new_n611_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n678_), .A2(new_n679_), .A3(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n576_), .A2(new_n517_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n627_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n686_), .A3(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n687_), .A2(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n691_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n685_), .A2(new_n686_), .A3(new_n693_), .A4(new_n689_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n631_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(G29gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n641_), .A2(new_n627_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n577_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n258_), .A2(new_n696_), .ZN(new_n699_));
  OAI22_X1  g498(.A1(new_n695_), .A2(new_n696_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT109), .ZN(G1328gat));
  INV_X1    g500(.A(new_n698_), .ZN(new_n702_));
  INV_X1    g501(.A(G36gat), .ZN(new_n703_));
  INV_X1    g502(.A(new_n482_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n702_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT45), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n482_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(new_n703_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n709_), .A2(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(KEYINPUT46), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n708_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n710_), .B1(new_n708_), .B2(new_n711_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1329gat));
  INV_X1    g513(.A(G43gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n702_), .A2(new_n715_), .A3(new_n428_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n429_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n715_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT47), .Z(G1330gat));
  NAND2_X1  g518(.A1(new_n692_), .A2(new_n694_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n464_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n722_), .A2(KEYINPUT111), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(KEYINPUT111), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(G50gat), .A3(new_n724_), .ZN(new_n725_));
  OR3_X1    g524(.A1(new_n698_), .A2(G50gat), .A3(new_n464_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1331gat));
  NAND2_X1  g526(.A1(new_n629_), .A2(new_n576_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n728_), .A2(KEYINPUT112), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(KEYINPUT112), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n483_), .A2(new_n516_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n729_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G57gat), .B1(new_n733_), .B2(new_n258_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n576_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n483_), .A2(new_n735_), .A3(new_n516_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n646_), .A2(new_n627_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n646_), .A2(KEYINPUT113), .A3(new_n627_), .A4(new_n736_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n258_), .A2(G57gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n734_), .B1(new_n741_), .B2(new_n742_), .ZN(G1332gat));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n733_), .A2(new_n744_), .A3(new_n704_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n741_), .A2(new_n704_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(G64gat), .ZN(new_n748_));
  AOI211_X1 g547(.A(KEYINPUT48), .B(new_n744_), .C1(new_n741_), .C2(new_n704_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1333gat));
  OR3_X1    g549(.A1(new_n732_), .A2(G71gat), .A3(new_n429_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n739_), .A2(new_n428_), .A3(new_n740_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G71gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G71gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(G1334gat));
  NAND3_X1  g557(.A1(new_n733_), .A2(new_n441_), .A3(new_n721_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n741_), .A2(new_n721_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(G78gat), .ZN(new_n762_));
  AOI211_X1 g561(.A(KEYINPUT50), .B(new_n441_), .C1(new_n741_), .C2(new_n721_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1335gat));
  NAND2_X1  g563(.A1(new_n736_), .A2(new_n697_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n258_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n735_), .A2(new_n627_), .A3(new_n516_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n685_), .A2(new_n768_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n258_), .A2(G85gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(G1336gat));
  AOI21_X1  g570(.A(G92gat), .B1(new_n766_), .B2(new_n704_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n704_), .A2(G92gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n769_), .B2(new_n773_), .ZN(G1337gat));
  NAND3_X1  g573(.A1(new_n766_), .A2(new_n529_), .A3(new_n428_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n769_), .A2(new_n428_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n776_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT115), .B1(new_n776_), .B2(G99gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g579(.A1(new_n685_), .A2(new_n721_), .A3(new_n768_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT116), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n685_), .A2(new_n783_), .A3(new_n768_), .A4(new_n721_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(G106gat), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT52), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n782_), .A2(new_n787_), .A3(G106gat), .A4(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n766_), .A2(new_n430_), .A3(new_n721_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1339gat));
  NOR2_X1   g594(.A1(new_n704_), .A2(new_n631_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n467_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n562_), .A2(KEYINPUT118), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n564_), .B2(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n561_), .A2(new_n555_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT55), .A3(new_n563_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n805_), .A2(KEYINPUT55), .A3(new_n563_), .A4(new_n802_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n568_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT56), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n807_), .A2(new_n811_), .A3(new_n568_), .A4(new_n808_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n810_), .A2(new_n516_), .A3(new_n570_), .A4(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n502_), .A2(new_n507_), .A3(new_n503_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n506_), .A2(new_n501_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n814_), .B(new_n512_), .C1(new_n507_), .C2(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n816_), .A2(new_n515_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n573_), .B2(new_n571_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n813_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n641_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n643_), .B1(new_n813_), .B2(new_n818_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT57), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n801_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n810_), .A2(new_n817_), .A3(new_n570_), .A4(new_n812_), .ZN(new_n826_));
  OR2_X1    g625(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n826_), .A2(new_n827_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n611_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n801_), .B1(new_n823_), .B2(KEYINPUT57), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n800_), .B1(new_n825_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n517_), .B2(new_n627_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n800_), .A2(KEYINPUT117), .A3(new_n516_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n612_), .B(new_n735_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT54), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n799_), .B1(new_n833_), .B2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G113gat), .B1(new_n839_), .B2(new_n516_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n833_), .A2(new_n838_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n798_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n830_), .A2(new_n822_), .A3(new_n824_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n800_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n838_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n842_), .A2(KEYINPUT59), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n516_), .A2(G113gat), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT121), .Z(new_n849_));
  AOI21_X1  g648(.A(new_n840_), .B1(new_n847_), .B2(new_n849_), .ZN(G1340gat));
  NAND2_X1  g649(.A1(new_n845_), .A2(new_n846_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n576_), .B(new_n851_), .C1(new_n839_), .C2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n735_), .B2(G120gat), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n839_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G120gat), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1341gat));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n842_), .B2(new_n800_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n800_), .A2(new_n860_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n851_), .B(new_n862_), .C1(new_n839_), .C2(new_n852_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT122), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n861_), .A2(new_n866_), .A3(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1342gat));
  INV_X1    g667(.A(new_n646_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G134gat), .B1(new_n839_), .B2(new_n869_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n611_), .A2(G134gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n847_), .B2(new_n871_), .ZN(G1343gat));
  AOI211_X1 g671(.A(new_n468_), .B(new_n797_), .C1(new_n833_), .C2(new_n838_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n516_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n576_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n627_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881_));
  AOI21_X1  g680(.A(G162gat), .B1(new_n873_), .B2(new_n869_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n468_), .B1(new_n833_), .B2(new_n838_), .ZN(new_n883_));
  INV_X1    g682(.A(G162gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n612_), .A2(new_n884_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n883_), .A2(new_n796_), .A3(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n881_), .B1(new_n882_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n796_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n884_), .B1(new_n888_), .B2(new_n646_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n873_), .A2(new_n885_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(KEYINPUT123), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n887_), .A2(new_n891_), .ZN(G1347gat));
  NAND2_X1  g691(.A1(new_n837_), .A2(KEYINPUT54), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n837_), .A2(KEYINPUT54), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n843_), .A2(new_n800_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n704_), .A2(new_n631_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n429_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n516_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT124), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n895_), .A2(new_n721_), .A3(new_n899_), .ZN(new_n900_));
  OR3_X1    g699(.A1(new_n900_), .A2(KEYINPUT125), .A3(new_n288_), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT125), .B1(new_n900_), .B2(new_n288_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n902_), .A3(KEYINPUT62), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n895_), .A2(new_n467_), .A3(new_n896_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n904_), .B(new_n516_), .C1(new_n270_), .C2(new_n269_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT125), .B(new_n906_), .C1(new_n900_), .C2(new_n288_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n903_), .A2(new_n905_), .A3(new_n907_), .ZN(G1348gat));
  AOI21_X1  g707(.A(new_n721_), .B1(new_n833_), .B2(new_n838_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n735_), .A2(new_n429_), .A3(new_n896_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n268_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n467_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n896_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n845_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n576_), .A2(new_n268_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  OR3_X1    g715(.A1(new_n911_), .A2(new_n916_), .A3(KEYINPUT126), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT126), .B1(new_n911_), .B2(new_n916_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1349gat));
  NOR3_X1   g718(.A1(new_n914_), .A2(new_n800_), .A3(new_n286_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n909_), .A2(new_n627_), .A3(new_n897_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n273_), .B2(new_n921_), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n904_), .A2(new_n282_), .A3(new_n869_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n904_), .A2(new_n611_), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n924_), .A2(KEYINPUT127), .A3(G190gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT127), .B1(new_n924_), .B2(G190gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n923_), .B1(new_n925_), .B2(new_n926_), .ZN(G1351gat));
  NAND2_X1  g726(.A1(new_n883_), .A2(new_n913_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n517_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n303_), .ZN(G1352gat));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n735_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(new_n306_), .ZN(G1353gat));
  INV_X1    g731(.A(new_n928_), .ZN(new_n933_));
  XOR2_X1   g732(.A(KEYINPUT63), .B(G211gat), .Z(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(new_n627_), .A3(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n928_), .B2(new_n800_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n935_), .A2(new_n937_), .ZN(G1354gat));
  AND3_X1   g737(.A1(new_n933_), .A2(G218gat), .A3(new_n611_), .ZN(new_n939_));
  AOI21_X1  g738(.A(G218gat), .B1(new_n933_), .B2(new_n869_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1355gat));
endmodule


