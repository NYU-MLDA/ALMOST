//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G71gat), .B(G78gat), .Z(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(KEYINPUT11), .B2(new_n204_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n207_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT9), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G85gat), .B(G92gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT9), .ZN(new_n224_));
  OR2_X1    g023(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n225_), .A2(KEYINPUT64), .A3(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT64), .B1(new_n225_), .B2(new_n226_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n221_), .B(new_n224_), .C1(new_n229_), .C2(G106gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n214_), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT65), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n213_), .A2(new_n215_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT7), .ZN(new_n237_));
  INV_X1    g036(.A(G99gat), .ZN(new_n238_));
  INV_X1    g037(.A(G106gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(new_n236_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n231_), .B1(new_n243_), .B2(new_n223_), .ZN(new_n244_));
  AOI211_X1 g043(.A(KEYINPUT8), .B(new_n222_), .C1(new_n242_), .C2(new_n216_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n230_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n211_), .A2(KEYINPUT12), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT66), .B(new_n230_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n210_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G230gat), .ZN(new_n252_));
  INV_X1    g051(.A(G233gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n245_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n240_), .A2(new_n241_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n259_), .B1(new_n216_), .B2(KEYINPUT65), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n222_), .B1(new_n260_), .B2(new_n236_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n258_), .B1(new_n261_), .B2(new_n231_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT66), .B1(new_n262_), .B2(new_n230_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n250_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n211_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT69), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n210_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269_));
  NOR3_X1   g068(.A1(new_n268_), .A2(new_n269_), .A3(KEYINPUT12), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n247_), .B(new_n257_), .C1(new_n267_), .C2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(new_n272_), .A3(new_n251_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n273_), .B(new_n254_), .C1(new_n272_), .C2(new_n251_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G120gat), .B(G148gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT5), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G176gat), .B(G204gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n271_), .A2(new_n274_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n203_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n282_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(KEYINPUT70), .A3(new_n280_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT13), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT71), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(KEYINPUT71), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n283_), .A2(new_n285_), .A3(KEYINPUT71), .A4(new_n287_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(KEYINPUT72), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT72), .B1(new_n290_), .B2(new_n291_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G8gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT78), .B(G8gat), .ZN(new_n298_));
  INV_X1    g097(.A(G1gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT14), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT79), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT80), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G15gat), .B(G22gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n303_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n297_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n305_), .A3(new_n296_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(G231gat), .A2(G233gat), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n312_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n211_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n210_), .A3(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G155gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT16), .ZN(new_n320_));
  XOR2_X1   g119(.A(G183gat), .B(G211gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT17), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n322_), .A2(new_n323_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT81), .B1(new_n318_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT81), .ZN(new_n328_));
  INV_X1    g127(.A(new_n326_), .ZN(new_n329_));
  AOI211_X1 g128(.A(new_n328_), .B(new_n329_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n325_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT82), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n325_), .B(KEYINPUT82), .C1(new_n327_), .C2(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G29gat), .B(G36gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT73), .ZN(new_n337_));
  XOR2_X1   g136(.A(G43gat), .B(G50gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT15), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT35), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G232gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT34), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n340_), .A2(new_n246_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n249_), .A2(new_n250_), .A3(new_n339_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n344_), .A2(new_n341_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n347_), .A2(new_n348_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G190gat), .B(G218gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(G134gat), .B(G162gat), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n352_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT36), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  OR3_X1    g156(.A1(new_n349_), .A2(new_n350_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n353_), .A2(new_n354_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT36), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT77), .B(KEYINPUT37), .Z(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(KEYINPUT76), .B(new_n360_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n358_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT37), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n335_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n295_), .A2(KEYINPUT83), .A3(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT24), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(G169gat), .B2(G176gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n374_), .B(KEYINPUT87), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n377_), .ZN(new_n381_));
  INV_X1    g180(.A(G183gat), .ZN(new_n382_));
  INV_X1    g181(.A(G190gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT23), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(G183gat), .A3(G190gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT25), .B(G183gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n379_), .A2(new_n381_), .A3(new_n387_), .A4(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G169gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n384_), .A2(KEYINPUT88), .A3(new_n386_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n395_), .B(KEYINPUT23), .C1(new_n382_), .C2(new_n383_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n393_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n391_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT89), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT89), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n391_), .A2(new_n402_), .A3(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405_));
  INV_X1    g204(.A(G43gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n404_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G127gat), .B(G134gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G113gat), .B(G120gat), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n410_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(KEYINPUT90), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n409_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n408_), .B(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G227gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(G15gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT30), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT31), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n417_), .A2(new_n422_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(G155gat), .A2(G162gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(KEYINPUT1), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(KEYINPUT1), .B2(new_n427_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G141gat), .A2(G148gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G141gat), .A2(G148gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(KEYINPUT2), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(KEYINPUT91), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT91), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n438_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT2), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n430_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n435_), .A2(new_n437_), .A3(new_n439_), .A4(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n426_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n443_), .A2(new_n427_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n434_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n416_), .A2(new_n446_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n429_), .A2(new_n433_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n411_), .A2(new_n412_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT4), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT4), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G225gat), .A2(G233gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n455_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT99), .B(G85gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT0), .B(G57gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n459_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n457_), .A2(new_n464_), .A3(new_n458_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n425_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G226gat), .A2(G233gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT19), .ZN(new_n471_));
  XOR2_X1   g270(.A(G197gat), .B(G204gat), .Z(new_n472_));
  OR2_X1    g271(.A1(new_n472_), .A2(KEYINPUT21), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(KEYINPUT21), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G211gat), .B(G218gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n474_), .A2(new_n475_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G169gat), .A2(G176gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n376_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n484_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n380_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n390_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n393_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n398_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n490_));
  OAI22_X1  g289(.A1(new_n488_), .A2(new_n397_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n482_), .B1(new_n491_), .B2(new_n478_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n471_), .B1(new_n480_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n401_), .A2(new_n479_), .A3(new_n403_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n471_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n496_), .B1(new_n491_), .B2(new_n478_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G8gat), .B(G36gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT18), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G64gat), .B(G92gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n494_), .A2(new_n497_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n471_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n403_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n402_), .B1(new_n391_), .B2(new_n399_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n478_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n491_), .A2(new_n478_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n471_), .A2(new_n496_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n507_), .A2(new_n503_), .A3(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n505_), .A2(KEYINPUT27), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT103), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT27), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n495_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n512_), .B1(new_n491_), .B2(new_n478_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n480_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n504_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n521_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n515_), .A2(new_n516_), .B1(new_n517_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n505_), .A2(KEYINPUT27), .A3(new_n514_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT103), .ZN(new_n525_));
  NOR2_X1   g324(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n253_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n446_), .A2(KEYINPUT29), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT94), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT94), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n530_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n448_), .A2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n529_), .B1(new_n479_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G78gat), .B(G106gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(KEYINPUT96), .Z(new_n543_));
  NAND3_X1  g342(.A1(new_n536_), .A2(new_n543_), .A3(new_n539_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n446_), .A2(KEYINPUT29), .ZN(new_n545_));
  XOR2_X1   g344(.A(G22gat), .B(G50gat), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n446_), .B2(KEYINPUT29), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n548_), .A2(new_n551_), .A3(new_n549_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n542_), .A2(new_n544_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n542_), .A2(KEYINPUT97), .A3(new_n544_), .A4(new_n555_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n543_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n540_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n544_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n555_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n558_), .A2(new_n559_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n523_), .A2(new_n525_), .A3(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n469_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n558_), .A2(new_n559_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n563_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n523_), .A2(new_n569_), .A3(new_n468_), .A4(new_n525_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n503_), .A2(KEYINPUT32), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n507_), .A2(new_n513_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT100), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT100), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n507_), .A2(new_n513_), .A3(new_n574_), .A4(new_n571_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT102), .ZN(new_n577_));
  INV_X1    g376(.A(new_n571_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n466_), .A2(new_n467_), .B1(new_n499_), .B2(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n576_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n577_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n464_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n582_), .A2(KEYINPUT33), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n456_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n447_), .A2(new_n450_), .A3(new_n456_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n464_), .ZN(new_n586_));
  OAI22_X1  g385(.A1(new_n582_), .A2(KEYINPUT33), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n583_), .A2(new_n587_), .A3(new_n522_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n580_), .A2(new_n581_), .A3(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n570_), .B1(new_n589_), .B2(new_n569_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n425_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n566_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n311_), .A2(new_n339_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT85), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n340_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT84), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n597_), .A2(new_n598_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n596_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n311_), .A2(new_n339_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n594_), .B1(new_n602_), .B2(new_n593_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G169gat), .B(G197gat), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n605_), .B(new_n606_), .Z(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n607_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n609_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(KEYINPUT86), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(KEYINPUT86), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n592_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n373_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n295_), .A2(new_n372_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT83), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n468_), .A2(G1gat), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n202_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n616_), .A2(KEYINPUT38), .A3(new_n619_), .A4(new_n621_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n611_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n293_), .A2(new_n294_), .A3(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n592_), .A2(new_n331_), .A3(new_n363_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n468_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n623_), .A2(new_n624_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT104), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n623_), .A2(new_n632_), .A3(new_n624_), .A4(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1324gat));
  NOR2_X1   g433(.A1(KEYINPUT106), .A2(KEYINPUT39), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n523_), .A2(new_n525_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n626_), .A2(new_n636_), .A3(new_n627_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(G8gat), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n637_), .B2(G8gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n635_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n641_), .ZN(new_n643_));
  XOR2_X1   g442(.A(KEYINPUT106), .B(KEYINPUT39), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n639_), .A3(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n616_), .A2(new_n298_), .A3(new_n619_), .A4(new_n636_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n642_), .A2(new_n645_), .A3(KEYINPUT40), .A4(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1325gat));
  XNOR2_X1  g450(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n628_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n419_), .B1(new_n654_), .B2(new_n425_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT108), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n655_), .A2(KEYINPUT108), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n653_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n658_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n652_), .A3(new_n656_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n425_), .A2(new_n419_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n659_), .B(new_n661_), .C1(new_n620_), .C2(new_n662_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n628_), .B2(new_n564_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n564_), .A2(G22gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n620_), .B2(new_n666_), .ZN(G1327gat));
  INV_X1    g466(.A(KEYINPUT110), .ZN(new_n668_));
  INV_X1    g467(.A(new_n335_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(new_n362_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n335_), .A2(KEYINPUT110), .A3(new_n363_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n672_), .A2(new_n295_), .A3(new_n615_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n468_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n365_), .A2(new_n370_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n592_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  INV_X1    g477(.A(new_n581_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n588_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n576_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n564_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n425_), .B1(new_n683_), .B2(new_n570_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n371_), .B(new_n678_), .C1(new_n684_), .C2(new_n566_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n677_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n626_), .A3(new_n335_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n686_), .A2(new_n626_), .A3(KEYINPUT44), .A4(new_n335_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n674_), .A2(G29gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n675_), .B1(new_n692_), .B2(new_n693_), .ZN(G1328gat));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n695_));
  INV_X1    g494(.A(new_n636_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n673_), .A2(new_n695_), .A3(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n672_), .A2(new_n295_), .A3(new_n615_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n697_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT45), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  AOI22_X1  g501(.A1(new_n698_), .A2(new_n701_), .B1(KEYINPUT111), .B2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n690_), .A2(new_n636_), .A3(new_n691_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G36gat), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n702_), .A2(KEYINPUT111), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n703_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  NAND4_X1  g508(.A1(new_n690_), .A2(G43gat), .A3(new_n425_), .A4(new_n691_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n406_), .B1(new_n699_), .B2(new_n591_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g512(.A(G50gat), .B1(new_n673_), .B2(new_n569_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n569_), .A2(G50gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n692_), .B2(new_n715_), .ZN(G1331gat));
  INV_X1    g515(.A(new_n592_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n625_), .ZN(new_n718_));
  NOR4_X1   g517(.A1(new_n295_), .A2(new_n718_), .A3(new_n335_), .A4(new_n371_), .ZN(new_n719_));
  INV_X1    g518(.A(G57gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n674_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n295_), .ZN(new_n722_));
  AND4_X1   g521(.A1(new_n669_), .A2(new_n717_), .A3(new_n362_), .A4(new_n614_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n722_), .A2(new_n674_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n720_), .B2(new_n724_), .ZN(G1332gat));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n719_), .A2(new_n726_), .A3(new_n636_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n723_), .A2(new_n722_), .A3(new_n636_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(G64gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G64gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n719_), .A2(new_n733_), .A3(new_n425_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n723_), .A2(new_n722_), .A3(new_n425_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G71gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G71gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1334gat));
  INV_X1    g538(.A(G78gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n719_), .A2(new_n740_), .A3(new_n569_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n723_), .A2(new_n722_), .A3(new_n569_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(G78gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(G78gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1335gat));
  NAND2_X1  g545(.A1(new_n335_), .A2(new_n625_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n294_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n292_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n686_), .A2(KEYINPUT112), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n686_), .A2(KEYINPUT112), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n468_), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n718_), .B(new_n295_), .C1(new_n671_), .C2(new_n670_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n218_), .A3(new_n674_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1336gat));
  AOI21_X1  g555(.A(G92gat), .B1(new_n754_), .B2(new_n636_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n752_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n636_), .A2(G92gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT113), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n757_), .B1(new_n758_), .B2(new_n760_), .ZN(G1337gat));
  OAI21_X1  g560(.A(G99gat), .B1(new_n752_), .B2(new_n591_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n591_), .A2(new_n229_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n754_), .A2(new_n763_), .B1(new_n764_), .B2(KEYINPUT51), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n764_), .A2(KEYINPUT51), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(G1338gat));
  NAND4_X1  g567(.A1(new_n686_), .A2(new_n749_), .A3(KEYINPUT115), .A4(new_n569_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G106gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n564_), .B1(new_n677_), .B2(new_n685_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT115), .B1(new_n771_), .B2(new_n749_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT52), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n749_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(G106gat), .A4(new_n769_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n773_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n754_), .A2(new_n239_), .A3(new_n569_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT53), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n779_), .A2(new_n783_), .A3(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1339gat));
  NOR3_X1   g584(.A1(new_n565_), .A2(new_n591_), .A3(new_n468_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n600_), .A2(new_n599_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n595_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n593_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n602_), .A2(new_n593_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n607_), .B1(new_n791_), .B2(new_n595_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n604_), .A2(new_n607_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n793_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n247_), .B(new_n251_), .C1(new_n267_), .C2(new_n270_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n254_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n247_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n265_), .A2(KEYINPUT69), .A3(new_n266_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n269_), .B1(new_n268_), .B2(KEYINPUT12), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT117), .B1(new_n800_), .B2(new_n257_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n796_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n271_), .A2(new_n804_), .A3(new_n802_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n278_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n797_), .B(new_n256_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT55), .B1(new_n810_), .B2(KEYINPUT117), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(new_n805_), .A3(new_n796_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n278_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n809_), .A2(KEYINPUT118), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n812_), .A2(new_n815_), .A3(KEYINPUT56), .A4(new_n278_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n281_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n794_), .B1(new_n814_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT57), .B1(new_n819_), .B2(new_n363_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(new_n817_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n271_), .A2(new_n804_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n823_), .A2(KEYINPUT55), .B1(new_n254_), .B2(new_n795_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n279_), .B1(new_n824_), .B2(new_n805_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n815_), .B1(new_n825_), .B2(KEYINPUT56), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n822_), .B1(new_n826_), .B2(new_n809_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n821_), .B(new_n362_), .C1(new_n827_), .C2(new_n794_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n820_), .A2(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n825_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n813_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n280_), .A4(new_n793_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT119), .B1(new_n825_), .B2(KEYINPUT56), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n807_), .A2(new_n831_), .A3(new_n808_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n836_), .A2(new_n837_), .B1(KEYINPUT56), .B2(new_n825_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n793_), .A2(new_n280_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n835_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n834_), .A2(new_n840_), .A3(new_n371_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n829_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n331_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n614_), .A2(new_n334_), .A3(new_n333_), .A4(new_n676_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n290_), .A2(new_n291_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n846_));
  OR3_X1    g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n787_), .B1(new_n843_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n611_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n669_), .B1(new_n829_), .B2(new_n841_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n853_), .A2(new_n849_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n787_), .A2(KEYINPUT59), .ZN(new_n855_));
  INV_X1    g654(.A(new_n331_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n829_), .B2(new_n841_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n786_), .B1(new_n857_), .B2(new_n849_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n854_), .A2(new_n855_), .B1(new_n858_), .B2(KEYINPUT59), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT120), .B(G113gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n612_), .A2(new_n613_), .A3(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT121), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n852_), .B1(new_n859_), .B2(new_n862_), .ZN(G1340gat));
  OAI21_X1  g662(.A(new_n855_), .B1(new_n853_), .B2(new_n849_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n851_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(G120gat), .B1(new_n866_), .B2(new_n295_), .ZN(new_n867_));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n295_), .B2(KEYINPUT60), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n851_), .B(new_n869_), .C1(KEYINPUT60), .C2(new_n868_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n867_), .A2(new_n870_), .ZN(G1341gat));
  INV_X1    g670(.A(G127gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n858_), .B2(new_n335_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(KEYINPUT122), .B(new_n872_), .C1(new_n858_), .C2(new_n335_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n331_), .A2(new_n872_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n875_), .A2(new_n876_), .B1(new_n859_), .B2(new_n877_), .ZN(G1342gat));
  AOI21_X1  g677(.A(G134gat), .B1(new_n851_), .B2(new_n363_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT123), .B(G134gat), .Z(new_n880_));
  NOR2_X1   g679(.A1(new_n676_), .A2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n859_), .B2(new_n881_), .ZN(G1343gat));
  AOI21_X1  g681(.A(new_n425_), .B1(new_n843_), .B2(new_n850_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n636_), .A2(new_n468_), .A3(new_n564_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n611_), .A3(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT124), .B(G141gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1344gat));
  NAND3_X1  g686(.A1(new_n883_), .A2(new_n722_), .A3(new_n884_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g688(.A1(new_n883_), .A2(new_n669_), .A3(new_n884_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  NAND3_X1  g691(.A1(new_n883_), .A2(new_n371_), .A3(new_n884_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G162gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n362_), .A2(G162gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n883_), .A2(new_n884_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1347gat));
  INV_X1    g696(.A(G169gat), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n636_), .A2(new_n468_), .A3(new_n564_), .A4(new_n425_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n611_), .B(new_n900_), .C1(new_n853_), .C2(new_n849_), .ZN(new_n901_));
  OAI211_X1 g700(.A(KEYINPUT62), .B(new_n898_), .C1(new_n901_), .C2(KEYINPUT22), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT62), .B1(new_n901_), .B2(KEYINPUT22), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n901_), .A2(KEYINPUT62), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n898_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n903_), .B1(new_n904_), .B2(new_n906_), .ZN(G1348gat));
  AND2_X1   g706(.A1(new_n854_), .A2(new_n900_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n722_), .ZN(new_n909_));
  INV_X1    g708(.A(G176gat), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n899_), .B1(new_n843_), .B2(new_n850_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n295_), .A2(new_n910_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n909_), .A2(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(G1349gat));
  AOI21_X1  g712(.A(G183gat), .B1(new_n911_), .B2(new_n669_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n331_), .A2(new_n388_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n908_), .B2(new_n915_), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n908_), .A2(new_n363_), .A3(new_n389_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n371_), .B(new_n900_), .C1(new_n853_), .C2(new_n849_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n918_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(KEYINPUT125), .B1(new_n918_), .B2(G190gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n917_), .B1(new_n919_), .B2(new_n920_), .ZN(G1351gat));
  NOR3_X1   g720(.A1(new_n696_), .A2(new_n674_), .A3(new_n564_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n883_), .A2(new_n611_), .A3(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT126), .B(G197gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1352gat));
  NAND3_X1  g724(.A1(new_n883_), .A2(new_n722_), .A3(new_n922_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G204gat), .ZN(G1353gat));
  OAI211_X1 g726(.A(new_n591_), .B(new_n922_), .C1(new_n857_), .C2(new_n849_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n856_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n931_), .A2(KEYINPUT127), .ZN(new_n932_));
  OR3_X1    g731(.A1(new_n928_), .A2(new_n930_), .A3(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n931_), .A2(KEYINPUT127), .ZN(new_n934_));
  OAI22_X1  g733(.A1(new_n928_), .A2(new_n930_), .B1(new_n934_), .B2(new_n932_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1354gat));
  OAI21_X1  g735(.A(G218gat), .B1(new_n928_), .B2(new_n676_), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n362_), .A2(G218gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n928_), .B2(new_n938_), .ZN(G1355gat));
endmodule


