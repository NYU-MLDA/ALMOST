//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(G169gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT80), .B(G183gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT23), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n209_), .B1(new_n211_), .B2(new_n216_), .ZN(new_n217_));
  OR3_X1    g016(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n208_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n218_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n210_), .A2(KEYINPUT25), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(KEYINPUT25), .B2(G183gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n222_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n215_), .B(KEYINPUT81), .ZN(new_n227_));
  INV_X1    g026(.A(new_n213_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n217_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(G15gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n230_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT31), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n230_), .B(new_n233_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT31), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n206_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT83), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n236_), .A2(new_n239_), .A3(new_n206_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT83), .B1(new_n245_), .B2(new_n240_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G127gat), .B(G134gat), .Z(new_n248_));
  XOR2_X1   g047(.A(G113gat), .B(G120gat), .Z(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n244_), .A2(new_n246_), .A3(new_n250_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT2), .ZN(new_n256_));
  INV_X1    g055(.A(G141gat), .ZN(new_n257_));
  INV_X1    g056(.A(G148gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n259_), .A2(new_n261_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT85), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n264_), .A2(KEYINPUT85), .A3(new_n268_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT29), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT84), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n267_), .B1(new_n266_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G141gat), .B(G148gat), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n273_), .A2(new_n274_), .A3(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G22gat), .B(G50gat), .Z(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n284_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n271_), .A2(new_n272_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(new_n274_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n255_), .B1(new_n285_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n283_), .A2(new_n284_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n255_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n274_), .A3(new_n286_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G78gat), .B(G106gat), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n295_), .A2(KEYINPUT91), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n295_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n289_), .A2(new_n298_), .A3(new_n293_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G211gat), .B(G218gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n301_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT21), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n302_), .A2(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT87), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G204gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G197gat), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n308_), .B(KEYINPUT21), .C1(new_n307_), .C2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(KEYINPUT88), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT21), .B1(new_n310_), .B2(new_n307_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(new_n307_), .B2(new_n305_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n306_), .B1(new_n312_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n302_), .A2(new_n303_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n318_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(G228gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n321_), .B(new_n323_), .C1(new_n274_), .C2(new_n287_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n311_), .A2(KEYINPUT88), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n314_), .A2(new_n315_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n319_), .B1(new_n327_), .B2(new_n306_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n273_), .A2(new_n282_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n324_), .B1(new_n323_), .B2(new_n331_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n297_), .A2(new_n299_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n332_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n250_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G225gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n287_), .A2(new_n251_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G85gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT0), .B(G57gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT96), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n337_), .A2(KEYINPUT4), .A3(new_n340_), .ZN(new_n348_));
  OR3_X1    g147(.A1(new_n287_), .A2(new_n251_), .A3(KEYINPUT4), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n338_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT96), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n341_), .A2(new_n351_), .A3(new_n345_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT97), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT97), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n347_), .A2(new_n355_), .A3(new_n350_), .A4(new_n352_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT33), .ZN(new_n357_));
  INV_X1    g156(.A(new_n345_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n338_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n339_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n354_), .A2(new_n356_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT18), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT93), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT20), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n373_), .B1(new_n328_), .B2(new_n230_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n209_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n227_), .A2(new_n228_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n225_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT25), .B(G183gat), .Z(new_n380_));
  OAI21_X1  g179(.A(new_n216_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n381_), .A2(new_n222_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n321_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n372_), .B1(new_n374_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT20), .B1(new_n321_), .B2(new_n383_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n370_), .B1(new_n328_), .B2(new_n230_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n367_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n317_), .A2(new_n230_), .A3(new_n320_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n378_), .A2(new_n382_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n390_), .B(KEYINPUT20), .C1(new_n328_), .C2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n371_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n370_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n230_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n321_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n373_), .B1(new_n328_), .B2(new_n391_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n366_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n389_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT94), .B(new_n367_), .C1(new_n385_), .C2(new_n388_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT95), .ZN(new_n404_));
  OR3_X1    g203(.A1(new_n361_), .A2(new_n404_), .A3(new_n357_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n404_), .B1(new_n361_), .B2(new_n357_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n362_), .A2(new_n403_), .A3(new_n405_), .A4(new_n406_), .ZN(new_n407_));
  OR3_X1    g206(.A1(new_n359_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n361_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n392_), .A2(new_n371_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n366_), .A2(KEYINPUT32), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n392_), .A2(new_n371_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT98), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n386_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n397_), .A2(KEYINPUT98), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n321_), .A2(new_n395_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n413_), .B1(new_n418_), .B2(new_n394_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n409_), .B(new_n412_), .C1(new_n419_), .C2(new_n411_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n336_), .B1(new_n407_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n401_), .A2(new_n422_), .A3(new_n402_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n410_), .B2(new_n366_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n419_), .B2(new_n366_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n426_), .A2(new_n335_), .A3(new_n409_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n254_), .B1(new_n421_), .B2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n335_), .A3(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT99), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n423_), .A2(new_n335_), .A3(new_n425_), .A4(KEYINPUT99), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n409_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n252_), .A2(new_n253_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n428_), .A2(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(G85gat), .A2(G92gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(G85gat), .A2(G92gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G99gat), .A2(G106gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT6), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(G99gat), .A3(G106gat), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G99gat), .A2(G106gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI22_X1  g247(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n440_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT8), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(KEYINPUT8), .B(new_n440_), .C1(new_n445_), .C2(new_n450_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT65), .B(G92gat), .Z(new_n455_));
  INV_X1    g254(.A(G85gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(KEYINPUT9), .ZN(new_n457_));
  AND2_X1   g256(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G106gat), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n455_), .A2(new_n457_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n440_), .A2(KEYINPUT9), .B1(new_n442_), .B2(new_n444_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n453_), .A2(new_n454_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT67), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n451_), .A2(new_n452_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT67), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n454_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G57gat), .B(G64gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G71gat), .B(G78gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT11), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(KEYINPUT11), .ZN(new_n473_));
  INV_X1    g272(.A(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n470_), .A2(KEYINPUT11), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT12), .B(new_n472_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n466_), .A2(new_n469_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT12), .ZN(new_n480_));
  INV_X1    g279(.A(new_n465_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n472_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G230gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT64), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n467_), .A2(new_n482_), .A3(new_n454_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n479_), .A2(new_n483_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n487_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n482_), .B1(new_n467_), .B2(new_n454_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n485_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G120gat), .B(G148gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT5), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G176gat), .B(G204gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n488_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n495_), .B(KEYINPUT68), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n498_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n499_));
  OR3_X1    g298(.A1(new_n497_), .A2(new_n499_), .A3(KEYINPUT13), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT13), .B1(new_n497_), .B2(new_n499_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G29gat), .B(G36gat), .Z(new_n503_));
  XOR2_X1   g302(.A(G43gat), .B(G50gat), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G29gat), .B(G36gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512_));
  INV_X1    g311(.A(G1gat), .ZN(new_n513_));
  INV_X1    g312(.A(G8gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G8gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n511_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n516_), .B(new_n517_), .Z(new_n520_));
  NAND3_X1  g319(.A1(new_n505_), .A2(KEYINPUT77), .A3(new_n508_), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT77), .B1(new_n505_), .B2(new_n508_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT78), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n519_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n521_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n518_), .B1(new_n528_), .B2(new_n522_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n525_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n527_), .A2(new_n530_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n534_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT79), .Z(new_n539_));
  AND3_X1   g338(.A1(new_n437_), .A2(new_n502_), .A3(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n541_));
  AND2_X1   g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT71), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n481_), .A2(new_n509_), .B1(new_n544_), .B2(new_n543_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n466_), .A2(new_n469_), .A3(new_n511_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n545_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n550_), .B1(KEYINPUT71), .B2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n548_), .A2(new_n549_), .A3(new_n546_), .A4(new_n545_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT72), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n554_), .A2(new_n555_), .A3(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n551_), .A2(KEYINPUT71), .ZN(new_n561_));
  AOI211_X1 g360(.A(new_n561_), .B(new_n547_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n553_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n559_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT72), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n558_), .B(KEYINPUT36), .Z(new_n567_));
  NAND3_X1  g366(.A1(new_n552_), .A2(new_n553_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(KEYINPUT73), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n566_), .A2(KEYINPUT73), .A3(KEYINPUT37), .A4(new_n568_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n518_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n482_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G127gat), .B(G155gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT17), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n583_), .A2(KEYINPUT17), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n578_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n584_), .B(KEYINPUT75), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n587_), .A2(KEYINPUT76), .A3(new_n577_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT76), .B1(new_n587_), .B2(new_n577_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n586_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n573_), .A2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n540_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n513_), .A3(new_n409_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT38), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n590_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n566_), .A2(new_n568_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n428_), .B2(new_n436_), .ZN(new_n599_));
  AND4_X1   g398(.A1(new_n596_), .A2(new_n599_), .A3(new_n502_), .A4(new_n538_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n513_), .B1(new_n600_), .B2(new_n409_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n594_), .B2(new_n593_), .ZN(G1324gat));
  NAND3_X1  g402(.A1(new_n592_), .A2(new_n514_), .A3(new_n426_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT100), .Z(new_n605_));
  AOI21_X1  g404(.A(new_n514_), .B1(new_n600_), .B2(new_n426_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT39), .Z(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(G1325gat));
  INV_X1    g409(.A(new_n254_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n232_), .B1(new_n600_), .B2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT41), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n592_), .A2(new_n232_), .A3(new_n611_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1326gat));
  INV_X1    g414(.A(G22gat), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n600_), .B2(new_n336_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT42), .Z(new_n618_));
  NAND3_X1  g417(.A1(new_n592_), .A2(new_n616_), .A3(new_n336_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1327gat));
  NOR2_X1   g419(.A1(new_n597_), .A2(new_n596_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n540_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(G29gat), .B1(new_n622_), .B2(new_n409_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n502_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n538_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n624_), .A2(new_n596_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n573_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(KEYINPUT43), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n437_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT103), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n437_), .A2(new_n631_), .A3(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n627_), .B1(new_n437_), .B2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n428_), .A2(new_n436_), .A3(KEYINPUT102), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n626_), .B1(new_n633_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT44), .B(new_n626_), .C1(new_n633_), .C2(new_n638_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n409_), .A2(G29gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n623_), .B1(new_n643_), .B2(new_n644_), .ZN(G1328gat));
  INV_X1    g444(.A(new_n622_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n426_), .ZN(new_n647_));
  OR3_X1    g446(.A1(new_n646_), .A2(G36gat), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT45), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n641_), .A2(new_n426_), .A3(new_n642_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(new_n651_), .A3(G36gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n650_), .B2(G36gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT46), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n649_), .B(KEYINPUT46), .C1(new_n652_), .C2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1329gat));
  NAND3_X1  g457(.A1(new_n643_), .A2(G43gat), .A3(new_n611_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n203_), .B1(new_n646_), .B2(new_n254_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g461(.A(G50gat), .B1(new_n622_), .B2(new_n336_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n336_), .A2(G50gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n643_), .B2(new_n664_), .ZN(G1331gat));
  AOI211_X1 g464(.A(new_n502_), .B(new_n538_), .C1(new_n428_), .C2(new_n436_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(new_n591_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G57gat), .B1(new_n667_), .B2(new_n409_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n539_), .A2(new_n590_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n599_), .A2(new_n624_), .A3(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n434_), .A2(KEYINPUT105), .ZN(new_n671_));
  MUX2_X1   g470(.A(KEYINPUT105), .B(new_n671_), .S(G57gat), .Z(new_n672_));
  AOI21_X1  g471(.A(new_n668_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT106), .Z(G1332gat));
  INV_X1    g473(.A(G64gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n670_), .B2(new_n426_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT48), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n667_), .A2(new_n675_), .A3(new_n426_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT107), .Z(G1333gat));
  INV_X1    g479(.A(G71gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n670_), .B2(new_n611_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT49), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n667_), .A2(new_n681_), .A3(new_n611_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1334gat));
  INV_X1    g484(.A(G78gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n670_), .B2(new_n336_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT50), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n667_), .A2(new_n686_), .A3(new_n336_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1335gat));
  NOR2_X1   g489(.A1(new_n633_), .A2(new_n638_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n624_), .A2(new_n590_), .A3(new_n625_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n456_), .B1(new_n693_), .B2(new_n409_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n666_), .A2(new_n621_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT108), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n434_), .A2(G85gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT109), .ZN(G1336gat));
  AOI21_X1  g498(.A(G92gat), .B1(new_n696_), .B2(new_n426_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n426_), .A2(new_n455_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n693_), .B2(new_n701_), .ZN(G1337gat));
  NAND2_X1  g501(.A1(new_n693_), .A2(new_n611_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n254_), .A2(new_n459_), .A3(new_n458_), .ZN(new_n704_));
  AOI22_X1  g503(.A1(new_n703_), .A2(G99gat), .B1(new_n696_), .B2(new_n704_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g505(.A(new_n461_), .B1(new_n693_), .B2(new_n336_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n707_), .A2(KEYINPUT52), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n696_), .A2(new_n461_), .A3(new_n336_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT110), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n696_), .A2(new_n711_), .A3(new_n461_), .A4(new_n336_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n707_), .A2(KEYINPUT52), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n708_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT53), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT53), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n708_), .A2(new_n713_), .A3(new_n717_), .A4(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1339gat));
  NAND3_X1  g518(.A1(new_n433_), .A2(new_n611_), .A3(new_n409_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n466_), .A2(new_n469_), .A3(new_n478_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n487_), .B1(new_n490_), .B2(KEYINPUT12), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n485_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(KEYINPUT55), .A3(new_n488_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n498_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n721_), .A2(new_n722_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT55), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n486_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n724_), .A2(new_n725_), .A3(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT56), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n498_), .A2(new_n730_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n724_), .A2(new_n728_), .A3(new_n732_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n497_), .B(new_n625_), .C1(new_n731_), .C2(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n497_), .A2(new_n499_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n526_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n519_), .A2(new_n524_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n524_), .A2(new_n529_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n526_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n740_), .B2(new_n534_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n736_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n742_), .A2(KEYINPUT112), .A3(new_n533_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n737_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n737_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n740_), .A2(new_n738_), .A3(new_n534_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT112), .B1(new_n742_), .B2(new_n533_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n535_), .B1(new_n750_), .B2(KEYINPUT113), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n735_), .A2(new_n746_), .A3(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n597_), .B1(new_n734_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT57), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT58), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n751_), .A2(new_n496_), .A3(new_n746_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(KEYINPUT114), .A2(new_n733_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n724_), .A2(new_n728_), .A3(new_n758_), .A4(new_n732_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n756_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n760_), .B2(KEYINPUT115), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n733_), .A2(KEYINPUT114), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n731_), .A2(new_n762_), .A3(new_n759_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n756_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT116), .B(new_n573_), .C1(new_n761_), .C2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n760_), .A2(KEYINPUT58), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n760_), .A2(KEYINPUT115), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n765_), .A2(new_n766_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n755_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT116), .B1(new_n773_), .B2(new_n573_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n754_), .B1(new_n770_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT117), .B(new_n754_), .C1(new_n770_), .C2(new_n774_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n590_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n669_), .B2(new_n502_), .ZN(new_n781_));
  NOR4_X1   g580(.A1(new_n539_), .A2(new_n624_), .A3(KEYINPUT111), .A4(new_n590_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n627_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n720_), .B1(new_n779_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n538_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n775_), .A2(new_n590_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n786_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n720_), .A2(KEYINPUT59), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT59), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n787_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n596_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n785_), .B1(new_n798_), .B2(new_n778_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT118), .B(KEYINPUT59), .C1(new_n799_), .C2(new_n720_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n794_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n801_), .A2(new_n539_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n789_), .B1(new_n802_), .B2(new_n788_), .ZN(G1340gat));
  INV_X1    g602(.A(G120gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n502_), .B2(KEYINPUT60), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n787_), .B(new_n805_), .C1(KEYINPUT60), .C2(new_n804_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n624_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n806_), .B1(new_n808_), .B2(new_n804_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT119), .B(new_n806_), .C1(new_n808_), .C2(new_n804_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(G1341gat));
  AOI21_X1  g612(.A(G127gat), .B1(new_n787_), .B2(new_n596_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n596_), .A2(G127gat), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT120), .Z(new_n816_));
  AOI21_X1  g615(.A(new_n814_), .B1(new_n801_), .B2(new_n816_), .ZN(G1342gat));
  AOI21_X1  g616(.A(G134gat), .B1(new_n787_), .B2(new_n598_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n573_), .A2(G134gat), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n819_), .B(KEYINPUT121), .Z(new_n820_));
  AOI21_X1  g619(.A(new_n818_), .B1(new_n801_), .B2(new_n820_), .ZN(G1343gat));
  NOR3_X1   g620(.A1(new_n799_), .A2(new_n611_), .A3(new_n335_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n409_), .A3(new_n647_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n625_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(new_n257_), .ZN(G1344gat));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n502_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(new_n258_), .ZN(G1345gat));
  NOR2_X1   g626(.A1(new_n823_), .A2(new_n590_), .ZN(new_n828_));
  XOR2_X1   g627(.A(KEYINPUT61), .B(G155gat), .Z(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1346gat));
  OAI21_X1  g629(.A(G162gat), .B1(new_n823_), .B2(new_n627_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n597_), .A2(G162gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n823_), .B2(new_n832_), .ZN(G1347gat));
  NOR2_X1   g632(.A1(new_n647_), .A2(new_n409_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n611_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n336_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n791_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G169gat), .B1(new_n837_), .B2(new_n625_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n838_), .A2(KEYINPUT62), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(KEYINPUT62), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT22), .B(G169gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n538_), .A2(new_n841_), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT122), .Z(new_n843_));
  OAI22_X1  g642(.A1(new_n839_), .A2(new_n840_), .B1(new_n837_), .B2(new_n843_), .ZN(G1348gat));
  INV_X1    g643(.A(new_n837_), .ZN(new_n845_));
  AOI21_X1  g644(.A(G176gat), .B1(new_n845_), .B2(new_n624_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(KEYINPUT123), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n799_), .A2(new_n336_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n835_), .A2(new_n219_), .A3(new_n502_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n847_), .A2(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(G1349gat));
  NAND3_X1  g650(.A1(new_n845_), .A2(new_n596_), .A3(new_n380_), .ZN(new_n852_));
  NOR4_X1   g651(.A1(new_n799_), .A2(new_n590_), .A3(new_n336_), .A4(new_n835_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n210_), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT124), .Z(G1350gat));
  OAI21_X1  g654(.A(G190gat), .B1(new_n837_), .B2(new_n627_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n598_), .A2(new_n225_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n837_), .B2(new_n857_), .ZN(G1351gat));
  NAND2_X1  g657(.A1(new_n822_), .A2(new_n834_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n625_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(G197gat), .Z(G1352gat));
  INV_X1    g660(.A(KEYINPUT126), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n859_), .B2(new_n502_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n862_), .B2(G204gat), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n822_), .A2(new_n624_), .A3(new_n834_), .A4(new_n865_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1353gat));
  NOR2_X1   g666(.A1(new_n859_), .A2(new_n590_), .ZN(new_n868_));
  OR2_X1    g667(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT63), .B(G211gat), .Z(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n868_), .B2(new_n871_), .ZN(G1354gat));
  OAI21_X1  g671(.A(G218gat), .B1(new_n859_), .B2(new_n627_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n597_), .A2(G218gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n822_), .A2(new_n834_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT127), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT127), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n873_), .A2(new_n878_), .A3(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1355gat));
endmodule


