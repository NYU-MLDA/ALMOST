//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT85), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(KEYINPUT1), .ZN(new_n206_));
  AND2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT82), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(new_n204_), .B2(KEYINPUT1), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT81), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT81), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G141gat), .A3(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(G141gat), .ZN(new_n217_));
  INV_X1    g016(.A(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n214_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n212_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT83), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n226_), .B1(new_n213_), .B2(KEYINPUT81), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n215_), .B1(new_n228_), .B2(KEYINPUT83), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n213_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n225_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n207_), .A2(new_n205_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n221_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT28), .B1(new_n235_), .B2(KEYINPUT29), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n227_), .A2(new_n228_), .B1(new_n230_), .B2(new_n213_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n233_), .B1(new_n237_), .B2(new_n225_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT28), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .A4(new_n221_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G22gat), .B(G50gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n236_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n242_), .B1(new_n236_), .B2(new_n241_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n203_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n245_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(KEYINPUT85), .A3(new_n243_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G197gat), .B(G204gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G211gat), .B(G218gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT84), .ZN(new_n251_));
  OAI211_X1 g050(.A(KEYINPUT21), .B(new_n249_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT21), .ZN(new_n253_));
  INV_X1    g052(.A(G218gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G211gat), .ZN(new_n255_));
  INV_X1    g054(.A(G211gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G218gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n253_), .B1(new_n258_), .B2(KEYINPUT84), .ZN(new_n259_));
  AND2_X1   g058(.A1(G197gat), .A2(G204gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G197gat), .A2(G204gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n250_), .B2(KEYINPUT21), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n252_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n265_), .B1(KEYINPUT29), .B2(new_n235_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G228gat), .A2(G233gat), .ZN(new_n267_));
  INV_X1    g066(.A(G78gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G106gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n266_), .B(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n246_), .A2(new_n248_), .A3(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT85), .B1(new_n247_), .B2(new_n243_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n272_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G127gat), .B(G134gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G113gat), .B(G120gat), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G113gat), .B(G120gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n235_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n238_), .A2(new_n284_), .A3(new_n221_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(KEYINPUT4), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G225gat), .A2(G233gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n284_), .B1(new_n238_), .B2(new_n221_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n238_), .A2(new_n284_), .A3(new_n221_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n293_), .A2(new_n290_), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n288_), .A2(new_n292_), .B1(new_n294_), .B2(new_n289_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G29gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G85gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT0), .B(G57gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n288_), .A2(new_n292_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n294_), .A2(new_n289_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n299_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G71gat), .B(G99gat), .ZN(new_n305_));
  INV_X1    g104(.A(G43gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT30), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(new_n285_), .ZN(new_n309_));
  XOR2_X1   g108(.A(KEYINPUT80), .B(KEYINPUT31), .Z(new_n310_));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT77), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(G169gat), .A3(G176gat), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n312_), .A2(new_n314_), .A3(KEYINPUT24), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(KEYINPUT76), .A2(G169gat), .A3(G176gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n315_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n312_), .A2(new_n314_), .A3(KEYINPUT24), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  INV_X1    g123(.A(G176gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n317_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT78), .B1(new_n322_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT25), .B(G183gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G190gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT24), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n327_), .A2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n321_), .A2(new_n328_), .A3(new_n336_), .A4(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n331_), .B(new_n332_), .C1(G183gat), .C2(G190gat), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n312_), .A2(new_n314_), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT22), .B(G169gat), .Z(new_n342_));
  OAI211_X1 g141(.A(new_n340_), .B(new_n341_), .C1(G176gat), .C2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT79), .B(G15gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G227gat), .A2(G233gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n339_), .A2(new_n343_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n310_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n310_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n348_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n309_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n309_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n300_), .B(new_n304_), .C1(new_n355_), .C2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n277_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n337_), .A2(KEYINPUT87), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT87), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT24), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n363_), .A2(new_n311_), .A3(new_n326_), .A4(new_n317_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n333_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n334_), .A2(new_n335_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n343_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n359_), .B1(new_n370_), .B2(new_n264_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n265_), .A2(new_n339_), .A3(new_n343_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n339_), .A2(new_n343_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n264_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n265_), .A2(new_n343_), .A3(new_n369_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n376_), .A2(new_n359_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .A4(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n370_), .B2(new_n264_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n259_), .A2(new_n263_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n339_), .A2(new_n343_), .B1(new_n385_), .B2(new_n252_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT88), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(G8gat), .B(G36gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT18), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n377_), .A2(new_n383_), .A3(new_n387_), .A4(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT27), .ZN(new_n393_));
  INV_X1    g192(.A(new_n391_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n376_), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n378_), .B2(new_n264_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n370_), .A2(KEYINPUT90), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n369_), .A2(new_n399_), .A3(new_n343_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n265_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n395_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n373_), .A2(new_n376_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n393_), .B1(new_n394_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n377_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n394_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT27), .B1(new_n408_), .B2(new_n392_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT92), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  AOI211_X1 g210(.A(KEYINPUT92), .B(KEYINPUT27), .C1(new_n408_), .C2(new_n392_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n358_), .B(new_n406_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n391_), .A2(KEYINPUT32), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n377_), .A2(new_n383_), .A3(new_n387_), .A4(new_n415_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n301_), .A2(new_n302_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n299_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n417_), .B(new_n418_), .C1(new_n421_), .C2(new_n303_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n294_), .A2(G225gat), .A3(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n288_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n289_), .B1(new_n286_), .B2(KEYINPUT4), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n423_), .B(new_n420_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n408_), .A2(new_n392_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n428_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n429_));
  AND4_X1   g228(.A1(new_n428_), .A2(new_n301_), .A3(new_n302_), .A4(new_n299_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n422_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n273_), .A2(new_n276_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT91), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT91), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n436_), .A3(new_n433_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n304_), .A2(new_n300_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n439_), .B(new_n406_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n355_), .A2(new_n356_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n414_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G120gat), .B(G148gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT5), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G176gat), .B(G204gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  INV_X1    g246(.A(KEYINPUT12), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(KEYINPUT68), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G57gat), .B(G64gat), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n452_));
  XOR2_X1   g251(.A(G71gat), .B(G78gat), .Z(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n452_), .A2(new_n453_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(KEYINPUT64), .B(G85gat), .Z(new_n457_));
  INV_X1    g256(.A(KEYINPUT9), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(G92gat), .ZN(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT10), .B(G99gat), .Z(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n270_), .ZN(new_n461_));
  OR2_X1    g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G85gat), .A2(G92gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(KEYINPUT9), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G99gat), .A3(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n459_), .A2(new_n461_), .A3(new_n464_), .A4(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT8), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT66), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT7), .ZN(new_n474_));
  INV_X1    g273(.A(G99gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n270_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT66), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n473_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G85gat), .B(G92gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT65), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n462_), .A2(new_n484_), .A3(new_n463_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n471_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n478_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n485_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT8), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n456_), .B(new_n470_), .C1(new_n487_), .C2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n479_), .A2(new_n469_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n486_), .A2(new_n471_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n478_), .B1(new_n469_), .B2(new_n472_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n489_), .B1(new_n495_), .B2(new_n480_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n496_), .B2(new_n471_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n456_), .B1(new_n497_), .B2(new_n470_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n449_), .B1(new_n492_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G230gat), .A2(G233gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n449_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n470_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n456_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n448_), .A2(KEYINPUT68), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n501_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n499_), .A2(new_n500_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n500_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n492_), .B2(new_n498_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT67), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT67), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n513_), .B(new_n510_), .C1(new_n492_), .C2(new_n498_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n447_), .B1(new_n509_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n447_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n508_), .A2(new_n512_), .A3(new_n514_), .A4(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT13), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(KEYINPUT13), .A3(new_n518_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524_));
  INV_X1    g323(.A(G1gat), .ZN(new_n525_));
  INV_X1    g324(.A(G8gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G1gat), .B(G8gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n456_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G127gat), .B(G155gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT17), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n538_), .A2(KEYINPUT17), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n533_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G29gat), .B(G36gat), .Z(new_n545_));
  XOR2_X1   g344(.A(G43gat), .B(G50gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT15), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n502_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n497_), .A2(new_n547_), .A3(new_n470_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT35), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n552_), .A2(KEYINPUT72), .A3(new_n553_), .A4(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT70), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n556_), .A2(new_n557_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n552_), .A2(KEYINPUT70), .A3(new_n553_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT71), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  AOI21_X1  g368(.A(new_n561_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n564_), .A2(new_n565_), .A3(new_n569_), .A4(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n565_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n569_), .A2(new_n565_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n562_), .A2(new_n563_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n573_), .B(new_n574_), .C1(new_n575_), .C2(new_n570_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(KEYINPUT73), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT37), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n572_), .A2(KEYINPUT73), .A3(new_n576_), .A4(KEYINPUT37), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n523_), .A2(new_n544_), .A3(new_n579_), .A4(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n530_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n547_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n548_), .A2(new_n530_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n548_), .A2(KEYINPUT75), .A3(new_n530_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n586_), .A2(G229gat), .A3(G233gat), .A4(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n549_), .A2(new_n530_), .A3(new_n551_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n583_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G113gat), .B(G141gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(G169gat), .B(G197gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n592_), .B(new_n595_), .Z(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n443_), .A2(new_n581_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT93), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n441_), .A2(new_n442_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n413_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n579_), .A2(new_n544_), .A3(new_n580_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n521_), .A2(new_n522_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n602_), .A2(new_n596_), .A3(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT93), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n202_), .B1(new_n600_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n598_), .A2(new_n599_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(KEYINPUT93), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(KEYINPUT94), .A3(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n608_), .A2(new_n525_), .A3(new_n438_), .A4(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n438_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n572_), .A2(new_n576_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n443_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n523_), .A2(new_n596_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n543_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n619_), .A2(KEYINPUT96), .A3(new_n621_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n616_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n525_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(KEYINPUT97), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n626_), .A2(new_n629_), .A3(new_n525_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n614_), .B(new_n615_), .C1(new_n628_), .C2(new_n630_), .ZN(G1324gat));
  INV_X1    g430(.A(KEYINPUT27), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n384_), .A2(new_n386_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n633_), .A2(new_n381_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n391_), .B1(new_n634_), .B2(new_n387_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n392_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT92), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n409_), .A2(new_n410_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n405_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G8gat), .B1(new_n622_), .B2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT39), .ZN(new_n642_));
  INV_X1    g441(.A(new_n640_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n608_), .A2(new_n526_), .A3(new_n643_), .A4(new_n611_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n642_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1325gat));
  NOR2_X1   g447(.A1(new_n600_), .A2(new_n607_), .ZN(new_n649_));
  INV_X1    g448(.A(G15gat), .ZN(new_n650_));
  INV_X1    g449(.A(new_n442_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n624_), .A2(new_n625_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n651_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(new_n654_), .B2(G15gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(G1326gat));
  INV_X1    g456(.A(G22gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n649_), .A2(new_n658_), .A3(new_n277_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n653_), .A2(new_n277_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(G22gat), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT42), .B(new_n658_), .C1(new_n653_), .C2(new_n277_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(G1327gat));
  NAND2_X1  g463(.A1(new_n618_), .A2(new_n543_), .ZN(new_n665_));
  NOR4_X1   g464(.A1(new_n443_), .A2(new_n597_), .A3(new_n604_), .A4(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n666_), .B2(new_n438_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n523_), .A2(new_n596_), .A3(new_n543_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n579_), .A2(new_n580_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n602_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n443_), .A2(new_n673_), .A3(KEYINPUT43), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT44), .B(new_n669_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT99), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n640_), .A2(new_n439_), .B1(new_n434_), .B2(KEYINPUT91), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n651_), .B1(new_n677_), .B2(new_n437_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n670_), .B(new_n671_), .C1(new_n678_), .C2(new_n414_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n443_), .B2(new_n673_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n668_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n676_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n681_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n438_), .A2(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n667_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(KEYINPUT46), .ZN(new_n692_));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n643_), .B1(new_n681_), .B2(KEYINPUT44), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n684_), .B2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n640_), .A2(G36gat), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT100), .B(KEYINPUT45), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT101), .Z(new_n699_));
  AND3_X1   g498(.A1(new_n666_), .A2(new_n697_), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n666_), .B2(new_n697_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n692_), .B1(new_n696_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n692_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n694_), .B1(new_n676_), .B2(new_n683_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n702_), .B(new_n705_), .C1(new_n706_), .C2(new_n693_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(G1329gat));
  NOR2_X1   g507(.A1(new_n442_), .A2(new_n306_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n679_), .A2(new_n680_), .ZN(new_n710_));
  AND4_X1   g509(.A1(new_n682_), .A2(new_n710_), .A3(KEYINPUT44), .A4(new_n669_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n682_), .B1(new_n681_), .B2(KEYINPUT44), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n687_), .B(new_n709_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n666_), .A2(new_n651_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n306_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n713_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1330gat));
  AOI21_X1  g518(.A(G50gat), .B1(new_n666_), .B2(new_n277_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n277_), .A2(G50gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n688_), .B2(new_n721_), .ZN(G1331gat));
  NOR2_X1   g521(.A1(new_n443_), .A2(new_n596_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n603_), .A2(new_n523_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT104), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n616_), .B1(new_n725_), .B2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G57gat), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n523_), .A2(new_n596_), .A3(new_n543_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n619_), .A2(G57gat), .A3(new_n438_), .A4(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT105), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT106), .ZN(G1332gat));
  INV_X1    g534(.A(G64gat), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n619_), .A2(new_n731_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n643_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT48), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n726_), .A2(new_n736_), .A3(new_n643_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1333gat));
  INV_X1    g540(.A(G71gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n737_), .B2(new_n651_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT49), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n726_), .A2(new_n742_), .A3(new_n651_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1334gat));
  AOI21_X1  g545(.A(new_n268_), .B1(new_n737_), .B2(new_n277_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT50), .Z(new_n748_));
  NAND3_X1  g547(.A1(new_n726_), .A2(new_n268_), .A3(new_n277_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1335gat));
  NOR4_X1   g549(.A1(new_n443_), .A2(new_n596_), .A3(new_n523_), .A4(new_n665_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n438_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n604_), .A2(new_n597_), .A3(new_n543_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n753_), .A2(new_n754_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n679_), .A2(new_n680_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n438_), .A2(new_n457_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n752_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT108), .ZN(G1336gat));
  AOI21_X1  g559(.A(G92gat), .B1(new_n751_), .B2(new_n643_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n643_), .A2(G92gat), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT109), .Z(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n757_), .B2(new_n763_), .ZN(G1337gat));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n765_), .A2(KEYINPUT51), .ZN(new_n766_));
  INV_X1    g565(.A(new_n757_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G99gat), .B1(new_n767_), .B2(new_n442_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n751_), .A2(new_n651_), .A3(new_n460_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n766_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n765_), .A2(KEYINPUT51), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n751_), .A2(new_n270_), .A3(new_n277_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n757_), .A2(new_n277_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(G106gat), .ZN(new_n776_));
  AOI211_X1 g575(.A(KEYINPUT52), .B(new_n270_), .C1(new_n757_), .C2(new_n277_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n773_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1339gat));
  NAND3_X1  g581(.A1(new_n640_), .A2(new_n651_), .A3(new_n438_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n596_), .A2(new_n518_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n501_), .B1(new_n504_), .B2(new_n491_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n449_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n510_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(KEYINPUT55), .A3(new_n508_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n499_), .A2(new_n507_), .A3(new_n790_), .A4(new_n500_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n789_), .A2(new_n447_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n517_), .A2(new_n793_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n789_), .A2(new_n791_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n785_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n588_), .A2(new_n591_), .A3(new_n595_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n586_), .A2(new_n590_), .A3(new_n587_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n590_), .B1(new_n582_), .B2(new_n547_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n595_), .B1(new_n589_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n798_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT57), .B(new_n617_), .C1(new_n797_), .C2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n796_), .A2(KEYINPUT115), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n789_), .A2(new_n810_), .A3(new_n791_), .A4(new_n795_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n794_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n518_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n805_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(new_n814_), .A3(KEYINPUT58), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n815_), .A2(new_n671_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT58), .B1(new_n812_), .B2(new_n814_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n808_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n617_), .B1(new_n797_), .B2(new_n806_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT113), .B(new_n617_), .C1(new_n797_), .C2(new_n806_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n544_), .B1(new_n819_), .B2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n605_), .A2(new_n597_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(KEYINPUT54), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n581_), .B2(new_n596_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n433_), .B(new_n784_), .C1(new_n826_), .C2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n815_), .A2(new_n671_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n807_), .B1(new_n837_), .B2(new_n817_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n543_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n832_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n841_), .A2(KEYINPUT59), .A3(new_n433_), .A4(new_n784_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n597_), .B1(new_n835_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(G113gat), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n596_), .A2(new_n844_), .ZN(new_n845_));
  OAI22_X1  g644(.A1(new_n843_), .A2(new_n844_), .B1(new_n833_), .B2(new_n845_), .ZN(G1340gat));
  AOI21_X1  g645(.A(new_n523_), .B1(new_n835_), .B2(new_n842_), .ZN(new_n847_));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n523_), .B2(KEYINPUT60), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(KEYINPUT60), .B2(new_n848_), .ZN(new_n850_));
  OAI22_X1  g649(.A1(new_n847_), .A2(new_n848_), .B1(new_n833_), .B2(new_n850_), .ZN(G1341gat));
  AOI21_X1  g650(.A(new_n543_), .B1(new_n835_), .B2(new_n842_), .ZN(new_n852_));
  INV_X1    g651(.A(G127gat), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n544_), .A2(new_n853_), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n852_), .A2(new_n853_), .B1(new_n833_), .B2(new_n854_), .ZN(G1342gat));
  NAND2_X1  g654(.A1(new_n835_), .A2(new_n842_), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT116), .B(G134gat), .Z(new_n857_));
  NOR2_X1   g656(.A1(new_n673_), .A2(new_n857_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n833_), .A2(new_n617_), .ZN(new_n859_));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n856_), .A2(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(G1343gat));
  NAND2_X1  g660(.A1(new_n816_), .A2(new_n818_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n825_), .A2(new_n862_), .A3(new_n807_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n832_), .B1(new_n863_), .B2(new_n543_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n277_), .A2(new_n442_), .A3(new_n438_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n864_), .A2(new_n643_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n596_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT117), .B(G141gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1344gat));
  NAND2_X1  g668(.A1(new_n866_), .A2(new_n604_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g670(.A1(new_n866_), .A2(new_n544_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  AOI21_X1  g673(.A(G162gat), .B1(new_n866_), .B2(new_n618_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n671_), .A2(G162gat), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(KEYINPUT118), .Z(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n866_), .B2(new_n877_), .ZN(G1347gat));
  OR2_X1    g677(.A1(new_n640_), .A2(new_n357_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT119), .Z(new_n880_));
  OAI211_X1 g679(.A(new_n433_), .B(new_n880_), .C1(new_n826_), .C2(new_n832_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G169gat), .B1(new_n881_), .B2(new_n597_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  OAI211_X1 g683(.A(KEYINPUT62), .B(G169gat), .C1(new_n881_), .C2(new_n597_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n881_), .A2(new_n597_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n884_), .B(new_n885_), .C1(new_n886_), .C2(new_n342_), .ZN(G1348gat));
  OAI21_X1  g686(.A(KEYINPUT120), .B1(new_n864_), .B2(new_n277_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n841_), .A2(new_n889_), .A3(new_n433_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n523_), .A2(new_n325_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n888_), .A2(new_n890_), .A3(new_n880_), .A4(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n325_), .B1(new_n881_), .B2(new_n523_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1349gat));
  NOR3_X1   g693(.A1(new_n881_), .A2(new_n334_), .A3(new_n543_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n888_), .A2(new_n890_), .A3(new_n544_), .A4(new_n880_), .ZN(new_n896_));
  INV_X1    g695(.A(G183gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n881_), .B2(new_n673_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n618_), .A2(new_n335_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n841_), .A2(new_n433_), .A3(new_n880_), .A4(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT121), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n899_), .A2(new_n905_), .A3(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1351gat));
  XNOR2_X1  g706(.A(KEYINPUT124), .B(G197gat), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n439_), .A2(new_n442_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n911_), .A2(KEYINPUT122), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(KEYINPUT122), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n912_), .A2(new_n643_), .A3(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n909_), .B1(new_n864_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n914_), .ZN(new_n916_));
  OAI211_X1 g715(.A(KEYINPUT123), .B(new_n916_), .C1(new_n826_), .C2(new_n832_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n908_), .B1(new_n918_), .B2(new_n596_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n908_), .ZN(new_n920_));
  AOI211_X1 g719(.A(new_n597_), .B(new_n920_), .C1(new_n915_), .C2(new_n917_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1352gat));
  NOR2_X1   g721(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n523_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n918_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  AOI211_X1 g726(.A(new_n927_), .B(new_n923_), .C1(new_n915_), .C2(new_n917_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1353gat));
  AND2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  NOR2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT126), .ZN(new_n933_));
  AOI211_X1 g732(.A(new_n930_), .B(new_n543_), .C1(new_n931_), .C2(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(KEYINPUT123), .B1(new_n841_), .B2(new_n916_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n917_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n934_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n933_), .A2(new_n931_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n918_), .B(new_n934_), .C1(new_n931_), .C2(new_n933_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1354gat));
  NAND3_X1  g740(.A1(new_n918_), .A2(new_n254_), .A3(new_n618_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n673_), .B1(new_n915_), .B2(new_n917_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n254_), .B2(new_n943_), .ZN(G1355gat));
endmodule


