//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_;
  INV_X1    g000(.A(KEYINPUT7), .ZN(new_n202_));
  INV_X1    g001(.A(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT6), .B1(new_n203_), .B2(new_n204_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  XOR2_X1   g013(.A(G85gat), .B(G92gat), .Z(new_n215_));
  AND3_X1   g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n215_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n207_), .A2(new_n218_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n205_), .A2(KEYINPUT66), .A3(new_n206_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n217_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n214_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n206_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n218_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(new_n212_), .A3(new_n220_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n215_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT67), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n216_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT65), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT64), .B(G85gat), .Z(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G92gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n232_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT10), .B(G99gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n212_), .B1(new_n237_), .B2(G106gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT68), .B1(new_n230_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n216_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n227_), .A2(new_n222_), .A3(new_n215_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT8), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n222_), .B1(new_n227_), .B2(new_n215_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n241_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n246_));
  INV_X1    g045(.A(new_n239_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n240_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G29gat), .B(G36gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G43gat), .B(G50gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(KEYINPUT70), .B(new_n241_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n229_), .A2(KEYINPUT8), .A3(new_n242_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT70), .B1(new_n256_), .B2(new_n241_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n247_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n252_), .B(KEYINPUT15), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G232gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT34), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n263_), .A2(KEYINPUT35), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n253_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT35), .A3(new_n263_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(KEYINPUT35), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n253_), .A2(new_n261_), .A3(new_n267_), .A4(new_n264_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G190gat), .B(G218gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(G134gat), .B(G162gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT36), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT74), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n266_), .A2(new_n268_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n266_), .A2(new_n268_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n271_), .B(KEYINPUT36), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT75), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n281_), .A3(new_n278_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n276_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT96), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT97), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290_));
  INV_X1    g089(.A(G169gat), .ZN(new_n291_));
  INV_X1    g090(.A(G176gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(KEYINPUT82), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(G169gat), .B2(G176gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n289_), .B1(new_n290_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT83), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT25), .B(G183gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT26), .B(G190gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(KEYINPUT81), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT24), .B1(new_n291_), .B2(new_n292_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n296_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n296_), .A2(new_n290_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n287_), .B(KEYINPUT23), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT83), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n302_), .A2(KEYINPUT81), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n299_), .A2(new_n306_), .A3(new_n310_), .A4(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(G169gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n287_), .A2(new_n288_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n287_), .A2(new_n288_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(G183gat), .B2(G190gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n314_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT88), .B(G197gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(G204gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT21), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n323_), .B1(G197gat), .B2(G204gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G197gat), .A2(G204gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n326_), .B1(new_n321_), .B2(G204gat), .ZN(new_n327_));
  OAI221_X1 g126(.A(new_n320_), .B1(new_n322_), .B2(new_n325_), .C1(KEYINPUT21), .C2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n320_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(KEYINPUT21), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n319_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT19), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n297_), .A2(new_n302_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n304_), .A2(KEYINPUT90), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n304_), .A2(KEYINPUT90), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n336_), .A2(new_n337_), .A3(new_n296_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n314_), .ZN(new_n339_));
  INV_X1    g138(.A(G183gat), .ZN(new_n340_));
  INV_X1    g139(.A(G190gat), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n289_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OAI22_X1  g141(.A1(new_n335_), .A2(new_n338_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT20), .B1(new_n343_), .B2(new_n331_), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n332_), .A2(new_n334_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n331_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n346_), .B(KEYINPUT20), .C1(new_n319_), .C2(new_n331_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n334_), .B2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G8gat), .B(G36gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT18), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n352_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n356_), .A2(KEYINPUT27), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n334_), .B1(new_n332_), .B2(new_n344_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n334_), .B2(new_n347_), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n352_), .B(KEYINPUT93), .Z(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n354_), .A2(new_n361_), .A3(KEYINPUT27), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT94), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n367_), .A2(KEYINPUT2), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(KEYINPUT2), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n368_), .A2(new_n371_), .A3(new_n372_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(KEYINPUT1), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n381_), .B(KEYINPUT85), .Z(new_n382_));
  INV_X1    g181(.A(new_n375_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT1), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n376_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AOI211_X1 g184(.A(new_n367_), .B(new_n369_), .C1(new_n382_), .C2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n387_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n380_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT29), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n331_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(G228gat), .A3(G233gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n331_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n366_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n396_), .A3(new_n366_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n391_), .A2(KEYINPUT29), .ZN(new_n401_));
  XOR2_X1   g200(.A(G22gat), .B(G50gat), .Z(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT28), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n401_), .B(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n397_), .B2(KEYINPUT89), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n398_), .A2(KEYINPUT89), .A3(new_n399_), .A4(new_n404_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G71gat), .B(G99gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G43gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G15gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n410_), .B(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n319_), .B(KEYINPUT30), .Z(new_n414_));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n414_), .A2(new_n415_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n413_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(new_n416_), .B2(new_n413_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G127gat), .B(G134gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G113gat), .B(G120gat), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(new_n421_), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT31), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n418_), .B(new_n423_), .C1(new_n416_), .C2(new_n413_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n380_), .A2(new_n390_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n422_), .B1(new_n430_), .B2(new_n388_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n422_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n389_), .A2(new_n432_), .A3(new_n380_), .A4(new_n390_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n433_), .A3(KEYINPUT91), .ZN(new_n434_));
  INV_X1    g233(.A(new_n430_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT91), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n432_), .A4(new_n389_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(KEYINPUT4), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n431_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n429_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n429_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G1gat), .B(G29gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(G85gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT0), .B(G57gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n441_), .A2(new_n443_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR4_X1   g251(.A1(new_n364_), .A2(new_n408_), .A3(new_n428_), .A4(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n408_), .A2(new_n454_), .A3(new_n357_), .A4(new_n363_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n352_), .A2(KEYINPUT32), .ZN(new_n456_));
  MUX2_X1   g255(.A(new_n359_), .B(new_n348_), .S(new_n456_), .Z(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT92), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n459_), .B1(new_n450_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n449_), .A2(KEYINPUT92), .A3(KEYINPUT33), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n434_), .A2(new_n437_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n447_), .B1(new_n464_), .B2(new_n442_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n438_), .A2(new_n440_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n465_), .B1(new_n466_), .B2(new_n442_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n356_), .B(new_n467_), .C1(new_n449_), .C2(KEYINPUT33), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n458_), .B1(new_n463_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n455_), .B1(new_n470_), .B2(new_n408_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n453_), .B1(new_n471_), .B2(new_n428_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n286_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G57gat), .B(G64gat), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n474_), .A2(KEYINPUT11), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(KEYINPUT11), .ZN(new_n476_));
  XOR2_X1   g275(.A(G71gat), .B(G78gat), .Z(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n476_), .A2(new_n477_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT69), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n240_), .A2(new_n248_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n483_));
  INV_X1    g282(.A(new_n480_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT12), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n482_), .A2(new_n483_), .B1(new_n258_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G230gat), .A2(G233gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n481_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n249_), .B2(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n246_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n490_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n482_), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n487_), .A2(new_n491_), .B1(new_n495_), .B2(new_n489_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G120gat), .B(G148gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT5), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G176gat), .B(G204gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT71), .B1(new_n496_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n482_), .A2(new_n483_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n258_), .A2(new_n486_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n503_), .A2(new_n488_), .A3(new_n504_), .A4(new_n494_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n495_), .A2(new_n489_), .ZN(new_n506_));
  AND4_X1   g305(.A1(KEYINPUT71), .A2(new_n505_), .A3(new_n506_), .A4(new_n501_), .ZN(new_n507_));
  OAI22_X1  g306(.A1(new_n502_), .A2(new_n507_), .B1(new_n496_), .B2(new_n501_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT13), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(KEYINPUT72), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(KEYINPUT72), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G1gat), .B(G8gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT76), .ZN(new_n514_));
  XOR2_X1   g313(.A(G15gat), .B(G22gat), .Z(new_n515_));
  NAND2_X1  g314(.A1(G1gat), .A2(G8gat), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(KEYINPUT14), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n514_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT77), .Z(new_n520_));
  XOR2_X1   g319(.A(new_n518_), .B(new_n520_), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(new_n480_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524_));
  XOR2_X1   g323(.A(G127gat), .B(G155gat), .Z(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT16), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G183gat), .B(G211gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n523_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(new_n484_), .B2(new_n521_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n528_), .B(new_n524_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n522_), .B2(new_n481_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n532_), .B1(new_n481_), .B2(new_n522_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n259_), .A2(new_n518_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n518_), .A2(new_n252_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n518_), .B(new_n252_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT80), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT79), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G169gat), .B(G197gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n544_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n512_), .A2(new_n534_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n473_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(G1gat), .B1(new_n553_), .B2(new_n454_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT38), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n512_), .A2(KEYINPUT73), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n510_), .A2(KEYINPUT73), .A3(new_n511_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n279_), .A2(KEYINPUT37), .A3(new_n275_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n283_), .B2(KEYINPUT37), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(new_n534_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT78), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n472_), .A2(new_n551_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n558_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(KEYINPUT95), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(KEYINPUT95), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n454_), .A2(G1gat), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n555_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n568_), .B2(new_n555_), .ZN(new_n571_));
  OAI221_X1 g370(.A(new_n554_), .B1(new_n555_), .B2(new_n568_), .C1(new_n570_), .C2(new_n571_), .ZN(G1324gat));
  INV_X1    g371(.A(G8gat), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n565_), .A2(new_n573_), .A3(new_n364_), .A4(new_n566_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT39), .ZN(new_n575_));
  INV_X1    g374(.A(new_n553_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n364_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n575_), .B1(new_n577_), .B2(G8gat), .ZN(new_n578_));
  AOI211_X1 g377(.A(KEYINPUT39), .B(new_n573_), .C1(new_n576_), .C2(new_n364_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n574_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n580_), .B(new_n582_), .ZN(G1325gat));
  OAI21_X1  g382(.A(G15gat), .B1(new_n553_), .B2(new_n428_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT41), .Z(new_n585_));
  INV_X1    g384(.A(G15gat), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n564_), .A2(new_n586_), .A3(new_n427_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(G1326gat));
  INV_X1    g387(.A(new_n408_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G22gat), .B1(new_n553_), .B2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT42), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n589_), .A2(G22gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT100), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n564_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(G1327gat));
  NAND2_X1  g394(.A1(new_n510_), .A2(new_n511_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n284_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n534_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n563_), .A2(new_n596_), .A3(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n454_), .A2(G29gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT103), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT44), .ZN(new_n604_));
  INV_X1    g403(.A(new_n560_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT43), .B1(new_n472_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT43), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n468_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n589_), .B1(new_n608_), .B2(new_n458_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n427_), .B1(new_n609_), .B2(new_n455_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n607_), .B(new_n560_), .C1(new_n610_), .C2(new_n453_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n512_), .A2(new_n551_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n614_), .A3(new_n534_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n613_), .B2(new_n534_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n604_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n534_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT101), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n620_), .A2(KEYINPUT44), .A3(new_n612_), .A4(new_n615_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n618_), .A2(new_n452_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n618_), .A2(KEYINPUT102), .A3(new_n452_), .A4(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G29gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n603_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT104), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n629_), .B(new_n603_), .C1(new_n624_), .C2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(G1328gat));
  NAND3_X1  g430(.A1(new_n618_), .A2(new_n364_), .A3(new_n621_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G36gat), .ZN(new_n633_));
  INV_X1    g432(.A(G36gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n600_), .A2(new_n634_), .A3(new_n364_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT45), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT46), .Z(G1329gat));
  AND2_X1   g437(.A1(new_n618_), .A2(new_n621_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(G43gat), .A3(new_n427_), .ZN(new_n640_));
  INV_X1    g439(.A(G43gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n600_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(new_n428_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g444(.A(G50gat), .B1(new_n600_), .B2(new_n408_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n408_), .A2(G50gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n639_), .B2(new_n647_), .ZN(G1331gat));
  NOR2_X1   g447(.A1(new_n472_), .A2(new_n550_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n512_), .A3(new_n562_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n452_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(G57gat), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n534_), .A2(new_n550_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n473_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n558_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n454_), .A2(new_n655_), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n654_), .A2(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(G1332gat));
  INV_X1    g459(.A(G64gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n658_), .B2(new_n364_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT48), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n651_), .A2(new_n661_), .A3(new_n364_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1333gat));
  INV_X1    g464(.A(KEYINPUT49), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n658_), .A2(new_n427_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(G71gat), .ZN(new_n668_));
  INV_X1    g467(.A(G71gat), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT49), .B(new_n669_), .C1(new_n658_), .C2(new_n427_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n427_), .A2(new_n669_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT106), .Z(new_n672_));
  OAI22_X1  g471(.A1(new_n668_), .A2(new_n670_), .B1(new_n650_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1334gat));
  INV_X1    g474(.A(G78gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n658_), .B2(new_n408_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT50), .Z(new_n678_));
  NAND3_X1  g477(.A1(new_n651_), .A2(new_n676_), .A3(new_n408_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1335gat));
  AND4_X1   g479(.A1(new_n512_), .A2(new_n612_), .A3(new_n534_), .A4(new_n551_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n233_), .A3(new_n452_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n558_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n683_), .A2(new_n599_), .A3(new_n649_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n452_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n686_), .B2(G85gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT108), .ZN(G1336gat));
  AOI21_X1  g487(.A(G92gat), .B1(new_n684_), .B2(new_n364_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n364_), .A2(G92gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT109), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n681_), .B2(new_n691_), .ZN(G1337gat));
  AOI21_X1  g491(.A(new_n203_), .B1(new_n681_), .B2(new_n427_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n428_), .A2(new_n237_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n684_), .B2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g495(.A1(new_n684_), .A2(new_n204_), .A3(new_n408_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT52), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n681_), .A2(new_n408_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(G106gat), .ZN(new_n700_));
  AOI211_X1 g499(.A(KEYINPUT52), .B(new_n204_), .C1(new_n681_), .C2(new_n408_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT53), .ZN(G1339gat));
  AND3_X1   g502(.A1(new_n605_), .A2(new_n509_), .A3(new_n656_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n550_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT111), .B(new_n550_), .C1(new_n502_), .C2(new_n507_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n503_), .A2(new_n494_), .A3(new_n504_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n489_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n487_), .A2(KEYINPUT55), .A3(new_n491_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT55), .B1(new_n487_), .B2(new_n491_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n715_), .B(new_n716_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT112), .B(KEYINPUT55), .C1(new_n487_), .C2(new_n491_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n500_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT113), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT56), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n713_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT114), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n713_), .B(new_n728_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n535_), .A2(new_n536_), .A3(new_n540_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n539_), .A2(new_n537_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n549_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n542_), .B2(new_n549_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n508_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n727_), .A2(new_n729_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n708_), .B1(new_n736_), .B2(new_n597_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT116), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT116), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n726_), .A2(KEYINPUT114), .B1(new_n508_), .B2(new_n734_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n284_), .B1(new_n740_), .B2(new_n729_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n741_), .B2(new_n708_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n736_), .A2(KEYINPUT57), .A3(new_n597_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n734_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n744_));
  AND2_X1   g543(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n745_));
  NOR2_X1   g544(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n721_), .B2(new_n746_), .ZN(new_n747_));
  OAI221_X1 g546(.A(new_n500_), .B1(KEYINPUT117), .B2(KEYINPUT56), .C1(new_n719_), .C2(new_n720_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n560_), .B1(new_n749_), .B2(KEYINPUT58), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT118), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(KEYINPUT58), .ZN(new_n753_));
  OAI211_X1 g552(.A(KEYINPUT118), .B(new_n560_), .C1(new_n749_), .C2(KEYINPUT58), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n738_), .A2(new_n742_), .A3(new_n743_), .A4(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n707_), .B1(new_n756_), .B2(new_n534_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n364_), .A2(new_n408_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n454_), .A2(new_n428_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT59), .B1(new_n757_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n743_), .A2(new_n755_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(new_n737_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n706_), .B1(new_n763_), .B2(new_n598_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT59), .ZN(new_n765_));
  INV_X1    g564(.A(new_n760_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n761_), .A2(new_n550_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G113gat), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT119), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n770_), .B1(new_n757_), .B2(new_n760_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n743_), .B(new_n755_), .C1(new_n737_), .C2(KEYINPUT116), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n741_), .A2(new_n739_), .A3(new_n708_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n534_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n706_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT119), .A3(new_n766_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n551_), .A2(G113gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n771_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n769_), .A2(new_n778_), .ZN(G1340gat));
  INV_X1    g578(.A(KEYINPUT60), .ZN(new_n780_));
  AOI21_X1  g579(.A(G120gat), .B1(new_n512_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n780_), .B2(G120gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n771_), .A2(new_n776_), .A3(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n761_), .A2(new_n683_), .A3(new_n767_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT120), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(G120gat), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n784_), .A2(KEYINPUT120), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(G1341gat));
  AOI21_X1  g587(.A(new_n760_), .B1(new_n774_), .B2(new_n706_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n598_), .B(new_n767_), .C1(new_n789_), .C2(new_n765_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G127gat), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n534_), .A2(G127gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n771_), .A2(new_n776_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n791_), .A2(KEYINPUT121), .A3(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1342gat));
  AND4_X1   g597(.A1(G134gat), .A2(new_n761_), .A3(new_n560_), .A4(new_n767_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n771_), .A2(new_n776_), .A3(new_n286_), .ZN(new_n800_));
  INV_X1    g599(.A(G134gat), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT122), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(KEYINPUT122), .A3(new_n801_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n799_), .B1(new_n804_), .B2(new_n805_), .ZN(G1343gat));
  NOR4_X1   g605(.A1(new_n364_), .A2(new_n589_), .A3(new_n454_), .A4(new_n427_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n757_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n550_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n683_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n809_), .B2(new_n598_), .ZN(new_n815_));
  NOR4_X1   g614(.A1(new_n757_), .A2(KEYINPUT123), .A3(new_n534_), .A4(new_n808_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT61), .B(G155gat), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n818_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n815_), .A2(new_n816_), .A3(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1346gat));
  INV_X1    g621(.A(G162gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n809_), .A2(new_n823_), .A3(new_n286_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n757_), .A2(new_n605_), .A3(new_n808_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1347gat));
  NAND2_X1  g627(.A1(new_n764_), .A2(new_n589_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n364_), .A2(new_n454_), .A3(new_n427_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(KEYINPUT22), .B(G169gat), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n550_), .A2(new_n832_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT125), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n831_), .A2(new_n550_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(G169gat), .ZN(new_n838_));
  AOI211_X1 g637(.A(KEYINPUT62), .B(new_n291_), .C1(new_n831_), .C2(new_n550_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n835_), .B1(new_n838_), .B2(new_n839_), .ZN(G1348gat));
  AOI21_X1  g639(.A(G176gat), .B1(new_n831_), .B2(new_n512_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n757_), .A2(new_n408_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n558_), .A2(new_n292_), .A3(new_n830_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(G1349gat));
  NOR2_X1   g643(.A1(new_n830_), .A2(new_n534_), .ZN(new_n845_));
  AOI21_X1  g644(.A(G183gat), .B1(new_n842_), .B2(new_n845_), .ZN(new_n846_));
  NOR4_X1   g645(.A1(new_n829_), .A2(new_n534_), .A3(new_n300_), .A4(new_n830_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1350gat));
  NAND2_X1  g647(.A1(new_n286_), .A2(new_n301_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT126), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n831_), .A2(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n829_), .A2(new_n605_), .A3(new_n830_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n341_), .ZN(G1351gat));
  NAND4_X1  g652(.A1(new_n364_), .A2(new_n454_), .A3(new_n408_), .A4(new_n428_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n757_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n550_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n683_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n598_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n861_));
  AND2_X1   g660(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n860_), .B2(new_n861_), .ZN(G1354gat));
  NAND2_X1  g663(.A1(new_n855_), .A2(new_n286_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT127), .B(G218gat), .Z(new_n866_));
  NOR2_X1   g665(.A1(new_n605_), .A2(new_n866_), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n865_), .A2(new_n866_), .B1(new_n855_), .B2(new_n867_), .ZN(G1355gat));
endmodule


