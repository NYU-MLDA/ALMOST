//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  OR3_X1    g007(.A1(new_n208_), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT25), .B1(new_n208_), .B2(KEYINPUT77), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n204_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n207_), .B1(new_n216_), .B2(KEYINPUT78), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n212_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT79), .B(G176gat), .Z(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT22), .B(G169gat), .ZN(new_n222_));
  AOI22_X1  g021(.A1(new_n221_), .A2(new_n222_), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n217_), .A2(new_n219_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT80), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G15gat), .B(G43gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT30), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n225_), .B(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G71gat), .B(G99gat), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G120gat), .ZN(new_n231_));
  INV_X1    g030(.A(G134gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G127gat), .ZN(new_n233_));
  INV_X1    g032(.A(G127gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G134gat), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n233_), .A2(new_n235_), .A3(KEYINPUT81), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT81), .B1(new_n233_), .B2(new_n235_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n236_), .A2(new_n237_), .A3(G113gat), .ZN(new_n238_));
  INV_X1    g037(.A(G113gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT81), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n234_), .A2(G134gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n232_), .A2(G127gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n233_), .A2(new_n235_), .A3(KEYINPUT81), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n239_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n231_), .B1(new_n238_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(G113gat), .B1(new_n236_), .B2(new_n237_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n239_), .A3(new_n244_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(G120gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT31), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  OR2_X1    g052(.A1(new_n230_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n230_), .A2(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT25), .B(G183gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n210_), .A2(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(new_n215_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n207_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n259_), .A2(new_n260_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n261_));
  INV_X1    g060(.A(G197gat), .ZN(new_n262_));
  INV_X1    g061(.A(G204gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT88), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT88), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G204gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n262_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G197gat), .A2(G204gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G211gat), .B(G218gat), .Z(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(KEYINPUT21), .A3(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n264_), .A2(new_n266_), .A3(new_n262_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT21), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(G197gat), .B2(G204gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n270_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT89), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n277_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n261_), .B(new_n271_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n271_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n280_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n283_), .B2(new_n278_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n281_), .B(KEYINPUT20), .C1(new_n284_), .C2(new_n224_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G226gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT19), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT90), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n281_), .A2(KEYINPUT20), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT90), .ZN(new_n290_));
  INV_X1    g089(.A(new_n287_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n217_), .A2(new_n219_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n220_), .A2(new_n223_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n271_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .A4(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT20), .B1(new_n284_), .B2(new_n261_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n294_), .A2(new_n295_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n287_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n288_), .A2(new_n297_), .A3(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G8gat), .B(G36gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT18), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G64gat), .ZN(new_n304_));
  INV_X1    g103(.A(G92gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n301_), .B(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n307_), .A2(KEYINPUT27), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n306_), .B(KEYINPUT96), .Z(new_n309_));
  OAI21_X1  g108(.A(new_n291_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n289_), .A2(new_n287_), .A3(new_n296_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n306_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n313_), .B(KEYINPUT27), .C1(new_n314_), .C2(new_n301_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n308_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT91), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n319_), .B1(new_n320_), .B2(KEYINPUT1), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(KEYINPUT82), .B(new_n319_), .C1(new_n320_), .C2(KEYINPUT1), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT83), .ZN(new_n325_));
  OR3_X1    g124(.A1(new_n319_), .A2(new_n325_), .A3(KEYINPUT1), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n319_), .B2(KEYINPUT1), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n323_), .A2(new_n324_), .A3(new_n326_), .A4(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(G141gat), .ZN(new_n330_));
  INV_X1    g129(.A(G148gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(new_n329_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT3), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT85), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n329_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT2), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n334_), .A2(new_n340_), .A3(new_n330_), .A4(new_n331_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n329_), .A2(new_n337_), .A3(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n336_), .A2(new_n339_), .A3(new_n341_), .A4(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n345_));
  XOR2_X1   g144(.A(G155gat), .B(G162gat), .Z(new_n346_));
  AND3_X1   g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n333_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n318_), .B1(new_n349_), .B2(new_n250_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n346_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT86), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n354_), .A2(new_n333_), .B1(new_n249_), .B2(new_n246_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n350_), .A2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n349_), .A2(new_n250_), .A3(KEYINPUT91), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT4), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n349_), .A2(new_n250_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n361_), .A2(KEYINPUT4), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT92), .ZN(new_n364_));
  INV_X1    g163(.A(new_n357_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n354_), .A2(new_n333_), .A3(new_n249_), .A4(new_n246_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n361_), .A3(new_n318_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n364_), .B1(new_n368_), .B2(new_n359_), .ZN(new_n369_));
  AOI211_X1 g168(.A(KEYINPUT92), .B(new_n360_), .C1(new_n365_), .C2(new_n367_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n363_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G1gat), .B(G29gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT0), .ZN(new_n373_));
  INV_X1    g172(.A(G57gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G85gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n363_), .B(new_n379_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n284_), .B1(KEYINPUT29), .B2(new_n349_), .ZN(new_n382_));
  INV_X1    g181(.A(G233gat), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n383_), .A2(KEYINPUT87), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(KEYINPUT87), .ZN(new_n385_));
  OAI21_X1  g184(.A(G228gat), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n382_), .B(new_n386_), .Z(new_n387_));
  OR2_X1    g186(.A1(new_n349_), .A2(KEYINPUT29), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G22gat), .B(G50gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT28), .ZN(new_n391_));
  XOR2_X1   g190(.A(G78gat), .B(G106gat), .Z(new_n392_));
  XOR2_X1   g191(.A(new_n391_), .B(new_n392_), .Z(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n389_), .B(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n317_), .A2(new_n381_), .A3(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n306_), .A2(KEYINPUT32), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n312_), .A2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n301_), .B2(new_n397_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n380_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT93), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT93), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n358_), .A2(new_n405_), .A3(new_n359_), .A4(new_n362_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n379_), .B1(new_n368_), .B2(new_n360_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n377_), .A2(new_n401_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n363_), .B(new_n409_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n402_), .A2(new_n408_), .A3(new_n307_), .A4(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n400_), .B1(new_n411_), .B2(KEYINPUT94), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n307_), .A2(new_n410_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT94), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n402_), .A4(new_n408_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n395_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n396_), .B1(new_n416_), .B2(KEYINPUT95), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT95), .ZN(new_n418_));
  AOI211_X1 g217(.A(new_n418_), .B(new_n395_), .C1(new_n412_), .C2(new_n415_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n256_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n395_), .A2(new_n316_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n256_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n381_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT97), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT97), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n421_), .A2(new_n425_), .A3(new_n381_), .A4(new_n422_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n420_), .A2(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT10), .B(G99gat), .Z(new_n429_));
  INV_X1    g228(.A(G106gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G85gat), .B(G92gat), .Z(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT9), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G99gat), .A2(G106gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OR3_X1    g237(.A1(new_n376_), .A2(new_n305_), .A3(KEYINPUT9), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n431_), .A2(new_n433_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT66), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT65), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  OR3_X1    g244(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n442_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n443_), .B(KEYINPUT65), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n449_), .A2(KEYINPUT66), .A3(new_n438_), .A4(new_n446_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n432_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n432_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT8), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT68), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n441_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(KEYINPUT68), .A3(new_n455_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G57gat), .B(G64gat), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n461_), .A2(KEYINPUT11), .ZN(new_n462_));
  XOR2_X1   g261(.A(G71gat), .B(G78gat), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(KEYINPUT11), .A3(new_n461_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(KEYINPUT11), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n462_), .A2(new_n466_), .A3(new_n463_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT12), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n460_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n456_), .A2(new_n440_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n468_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n456_), .A2(new_n440_), .A3(new_n468_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n474_), .B1(new_n475_), .B2(new_n469_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G230gat), .A2(G233gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n477_), .B(KEYINPUT64), .Z(new_n478_));
  NAND3_X1  g277(.A1(new_n471_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n474_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n480_), .B1(new_n481_), .B2(new_n475_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n483_));
  XNOR2_X1  g282(.A(G120gat), .B(G148gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G176gat), .B(G204gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  NAND3_X1  g286(.A1(new_n479_), .A2(new_n482_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT70), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n492_), .A2(KEYINPUT13), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(KEYINPUT13), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G29gat), .B(G36gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G43gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT71), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n499_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(G50gat), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(G50gat), .B1(new_n500_), .B2(new_n501_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506_));
  INV_X1    g305(.A(G1gat), .ZN(new_n507_));
  INV_X1    g306(.A(G8gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT14), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G1gat), .B(G8gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G229gat), .A2(G233gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n498_), .B(new_n499_), .ZN(new_n521_));
  INV_X1    g320(.A(G50gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT72), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n502_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n524_), .B1(new_n523_), .B2(new_n502_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n520_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT72), .B1(new_n503_), .B2(new_n504_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(KEYINPUT15), .A3(new_n525_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n512_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n513_), .A2(new_n517_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n519_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G113gat), .B(G141gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G169gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(new_n262_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n529_), .A2(KEYINPUT15), .A3(new_n525_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT15), .B1(new_n529_), .B2(new_n525_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n514_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n532_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(new_n519_), .A3(new_n536_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n538_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n496_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT34), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n528_), .A2(new_n530_), .B1(new_n459_), .B2(new_n458_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n472_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n505_), .A2(new_n553_), .B1(new_n550_), .B2(new_n549_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n551_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(KEYINPUT36), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n460_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n551_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n554_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n556_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n559_), .B(KEYINPUT36), .Z(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT73), .Z(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n556_), .B2(new_n563_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT37), .B1(new_n565_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n556_), .A2(new_n563_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n566_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n564_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n512_), .B(KEYINPUT75), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n473_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n580_));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n578_), .B1(new_n579_), .B2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(KEYINPUT17), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n585_), .B1(new_n586_), .B2(new_n578_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n574_), .A2(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n428_), .A2(new_n546_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n381_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n507_), .A3(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT38), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n571_), .A2(new_n564_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n428_), .A2(KEYINPUT98), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT98), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n420_), .A2(new_n427_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n597_), .B2(new_n593_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n587_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n546_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n590_), .A3(new_n601_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n602_), .A2(KEYINPUT99), .A3(G1gat), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT99), .B1(new_n602_), .B2(G1gat), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n592_), .B1(new_n603_), .B2(new_n604_), .ZN(G1324gat));
  NAND3_X1  g404(.A1(new_n589_), .A2(new_n508_), .A3(new_n316_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n316_), .B(new_n601_), .C1(new_n595_), .C2(new_n598_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n607_), .A2(new_n608_), .A3(G8gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n607_), .B2(G8gat), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n606_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(G1325gat));
  NAND3_X1  g412(.A1(new_n599_), .A2(new_n422_), .A3(new_n601_), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(G15gat), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(G15gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n589_), .A2(new_n617_), .A3(new_n422_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n615_), .B1(new_n614_), .B2(G15gat), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1326gat));
  INV_X1    g420(.A(G22gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n589_), .A2(new_n622_), .A3(new_n395_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n599_), .A2(new_n395_), .A3(new_n601_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G22gat), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(KEYINPUT42), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(KEYINPUT42), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(G1327gat));
  NAND3_X1  g427(.A1(new_n496_), .A2(new_n600_), .A3(new_n545_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n428_), .A2(new_n593_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G29gat), .B1(new_n630_), .B2(new_n590_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n574_), .B(KEYINPUT102), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n597_), .B2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n574_), .A2(KEYINPUT43), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n420_), .B2(new_n427_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n629_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT44), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n640_), .A2(G29gat), .A3(new_n590_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n639_), .A2(KEYINPUT44), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n631_), .B1(new_n641_), .B2(new_n642_), .ZN(G1328gat));
  INV_X1    g442(.A(KEYINPUT46), .ZN(new_n644_));
  INV_X1    g443(.A(G36gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n317_), .B1(new_n639_), .B2(KEYINPUT44), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n642_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n630_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n316_), .A2(new_n645_), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n648_), .A2(KEYINPUT45), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT45), .B1(new_n648_), .B2(new_n649_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT103), .B(new_n644_), .C1(new_n647_), .C2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n640_), .A2(new_n316_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n639_), .A2(KEYINPUT44), .ZN(new_n655_));
  OAI21_X1  g454(.A(G36gat), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n650_), .A2(new_n651_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n644_), .A2(KEYINPUT103), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n653_), .A2(new_n659_), .ZN(G1329gat));
  INV_X1    g459(.A(G43gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(new_n648_), .B2(new_n256_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n640_), .A2(G43gat), .A3(new_n422_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(new_n655_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT47), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n666_), .B(new_n662_), .C1(new_n663_), .C2(new_n655_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1330gat));
  AOI21_X1  g467(.A(G50gat), .B1(new_n630_), .B2(new_n395_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n395_), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n522_), .B(new_n670_), .C1(new_n639_), .C2(KEYINPUT44), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n671_), .B2(new_n642_), .ZN(G1331gat));
  INV_X1    g471(.A(new_n545_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n495_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n600_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n599_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G57gat), .B1(new_n676_), .B2(new_n381_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n428_), .A2(new_n588_), .A3(new_n674_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n678_), .A2(new_n374_), .A3(new_n590_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1332gat));
  INV_X1    g479(.A(G64gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(new_n681_), .A3(new_n316_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G64gat), .B1(new_n676_), .B2(new_n317_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT48), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(KEYINPUT48), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n682_), .B1(new_n684_), .B2(new_n685_), .ZN(G1333gat));
  INV_X1    g485(.A(G71gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n678_), .A2(new_n687_), .A3(new_n422_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G71gat), .B1(new_n676_), .B2(new_n256_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(KEYINPUT49), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(KEYINPUT49), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(G1334gat));
  INV_X1    g491(.A(G78gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n678_), .A2(new_n693_), .A3(new_n395_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G78gat), .B1(new_n676_), .B2(new_n670_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT50), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT50), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(G1335gat));
  NOR2_X1   g497(.A1(new_n674_), .A2(new_n587_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n597_), .A2(new_n594_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G85gat), .B1(new_n701_), .B2(new_n590_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n633_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n420_), .B2(new_n427_), .ZN(new_n704_));
  OAI22_X1  g503(.A1(new_n428_), .A2(new_n636_), .B1(new_n704_), .B2(new_n632_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n699_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n590_), .A2(G85gat), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT104), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n702_), .B1(new_n706_), .B2(new_n708_), .ZN(G1336gat));
  NAND3_X1  g508(.A1(new_n701_), .A2(new_n305_), .A3(new_n316_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n706_), .A2(new_n316_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n305_), .ZN(G1337gat));
  NAND3_X1  g511(.A1(new_n701_), .A2(new_n429_), .A3(new_n422_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n706_), .A2(new_n422_), .ZN(new_n714_));
  INV_X1    g513(.A(G99gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n713_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g516(.A(KEYINPUT107), .B(KEYINPUT53), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n395_), .B(new_n699_), .C1(new_n634_), .C2(new_n637_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT106), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n705_), .A2(new_n721_), .A3(new_n395_), .A4(new_n699_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(G106gat), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n720_), .A2(KEYINPUT52), .A3(new_n722_), .A4(G106gat), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n670_), .A2(G106gat), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n700_), .A2(KEYINPUT105), .A3(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT105), .B1(new_n700_), .B2(new_n728_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  AND4_X1   g530(.A1(new_n718_), .A2(new_n725_), .A3(new_n726_), .A4(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n731_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n718_), .B1(new_n734_), .B2(new_n726_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n732_), .A2(new_n735_), .ZN(G1339gat));
  OR3_X1    g535(.A1(new_n495_), .A2(new_n588_), .A3(new_n545_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT108), .B(KEYINPUT54), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OR3_X1    g539(.A1(new_n737_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n740_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n737_), .B2(new_n740_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT57), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n536_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n513_), .A2(new_n518_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n531_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n544_), .A2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n492_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n479_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n471_), .A2(new_n476_), .A3(KEYINPUT55), .A4(new_n478_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n471_), .A2(new_n476_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n480_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n753_), .A3(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n487_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n752_), .A2(new_n755_), .A3(KEYINPUT111), .A4(new_n753_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(KEYINPUT56), .A3(new_n759_), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT112), .B(KEYINPUT56), .C1(new_n758_), .C2(new_n759_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n756_), .A2(new_n757_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n487_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n759_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n760_), .B1(new_n761_), .B2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n533_), .A2(new_n537_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n536_), .B1(new_n543_), .B2(new_n519_), .ZN(new_n770_));
  OAI211_X1 g569(.A(KEYINPUT110), .B(new_n488_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT110), .B1(new_n545_), .B2(new_n488_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n750_), .B1(new_n768_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n745_), .B1(new_n775_), .B2(new_n594_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n544_), .A2(new_n488_), .A3(new_n748_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n758_), .A2(KEYINPUT56), .A3(new_n759_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n758_), .B2(new_n759_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n778_), .B(KEYINPUT58), .C1(new_n779_), .C2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n574_), .B1(new_n781_), .B2(KEYINPUT114), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n765_), .A2(new_n766_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n777_), .B1(new_n783_), .B2(new_n760_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(KEYINPUT58), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n784_), .A2(KEYINPUT113), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n784_), .B2(KEYINPUT113), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n782_), .B(new_n786_), .C1(new_n787_), .C2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n776_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n768_), .A2(new_n774_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n492_), .A2(new_n749_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT57), .A3(new_n593_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT115), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n775_), .A2(new_n594_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(KEYINPUT57), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n791_), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n600_), .B1(new_n800_), .B2(KEYINPUT116), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n776_), .A2(new_n790_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n798_), .B1(new_n797_), .B2(KEYINPUT57), .ZN(new_n803_));
  NOR4_X1   g602(.A1(new_n775_), .A2(KEYINPUT115), .A3(new_n745_), .A4(new_n594_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n802_), .B(KEYINPUT116), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n744_), .B1(new_n801_), .B2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n421_), .A2(new_n590_), .A3(new_n422_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n239_), .B1(new_n810_), .B2(new_n673_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT117), .B(new_n239_), .C1(new_n810_), .C2(new_n673_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n744_), .B1(new_n587_), .B2(new_n800_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n809_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n821_));
  XOR2_X1   g620(.A(KEYINPUT119), .B(G113gat), .Z(new_n822_));
  NOR2_X1   g621(.A1(new_n673_), .A2(new_n822_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n813_), .A2(new_n814_), .B1(new_n821_), .B2(new_n823_), .ZN(G1340gat));
  NAND2_X1  g623(.A1(new_n817_), .A2(new_n820_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n495_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT120), .B1(new_n816_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n496_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n600_), .A3(new_n805_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n808_), .B1(new_n833_), .B2(new_n744_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n828_), .B(new_n829_), .C1(new_n834_), .C2(new_n815_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n827_), .A2(G120gat), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n496_), .B2(G120gat), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n834_), .B(new_n838_), .C1(new_n837_), .C2(G120gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(G1341gat));
  NAND2_X1  g639(.A1(new_n810_), .A2(KEYINPUT59), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(new_n587_), .A3(new_n825_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G127gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n834_), .A2(new_n234_), .A3(new_n587_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1342gat));
  INV_X1    g644(.A(new_n574_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n841_), .A2(new_n846_), .A3(new_n825_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G134gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n834_), .A2(new_n232_), .A3(new_n594_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1343gat));
  INV_X1    g649(.A(new_n807_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n670_), .A2(new_n422_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n590_), .A3(new_n317_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n851_), .A2(new_n673_), .A3(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(new_n330_), .ZN(G1344gat));
  NOR3_X1   g654(.A1(new_n851_), .A2(new_n496_), .A3(new_n853_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT121), .B(G148gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n856_), .B(new_n858_), .ZN(G1345gat));
  NOR3_X1   g658(.A1(new_n851_), .A2(new_n600_), .A3(new_n853_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT122), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n860_), .B(new_n863_), .ZN(G1346gat));
  NOR2_X1   g663(.A1(new_n851_), .A2(new_n853_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G162gat), .B1(new_n865_), .B2(new_n594_), .ZN(new_n866_));
  INV_X1    g665(.A(G162gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n703_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n865_), .B2(new_n868_), .ZN(G1347gat));
  INV_X1    g668(.A(G169gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n317_), .A2(new_n590_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n422_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n545_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT123), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n395_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n870_), .B1(new_n817_), .B2(new_n876_), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT62), .Z(new_n878_));
  NAND3_X1  g677(.A1(new_n817_), .A2(new_n670_), .A3(new_n873_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n545_), .A2(new_n222_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT124), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n878_), .B1(new_n879_), .B2(new_n881_), .ZN(G1348gat));
  OR2_X1    g681(.A1(new_n879_), .A2(new_n496_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n851_), .A2(new_n395_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n873_), .A2(new_n495_), .A3(G176gat), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n221_), .A2(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1349gat));
  NOR3_X1   g685(.A1(new_n872_), .A2(new_n257_), .A3(new_n600_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n817_), .A2(new_n670_), .A3(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT125), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n884_), .A2(new_n587_), .A3(new_n873_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n208_), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n879_), .B2(new_n574_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n594_), .A2(new_n210_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n879_), .B2(new_n893_), .ZN(G1351gat));
  NAND2_X1  g693(.A1(new_n852_), .A2(new_n871_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n833_), .B2(new_n744_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n545_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g697(.A1(new_n264_), .A2(new_n266_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n896_), .A2(new_n900_), .A3(new_n495_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n896_), .A2(KEYINPUT127), .A3(new_n900_), .A4(new_n495_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n807_), .A2(new_n852_), .A3(new_n871_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n496_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n896_), .A2(KEYINPUT126), .A3(new_n495_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(G204gat), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n905_), .A2(new_n910_), .ZN(G1353gat));
  OR2_X1    g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  AND4_X1   g712(.A1(new_n587_), .A2(new_n896_), .A3(new_n912_), .A4(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n896_), .B2(new_n587_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1354gat));
  OR3_X1    g715(.A1(new_n907_), .A2(G218gat), .A3(new_n593_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G218gat), .B1(new_n907_), .B2(new_n574_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1355gat));
endmodule


