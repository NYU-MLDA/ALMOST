//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n923_, new_n924_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G1gat), .B(G8gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT75), .ZN(new_n205_));
  INV_X1    g004(.A(G15gat), .ZN(new_n206_));
  INV_X1    g005(.A(G22gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G15gat), .A2(G22gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G1gat), .A2(G8gat), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n208_), .A2(new_n209_), .B1(KEYINPUT14), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n205_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G43gat), .B(G50gat), .Z(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n212_), .A2(new_n219_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n203_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n212_), .A2(new_n219_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT70), .B(KEYINPUT15), .Z(new_n224_));
  XNOR2_X1  g023(.A(new_n219_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n205_), .A2(new_n211_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n205_), .A2(new_n211_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n223_), .A2(new_n228_), .A3(new_n202_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n222_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G113gat), .B(G141gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G169gat), .B(G197gat), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n231_), .B(new_n232_), .Z(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT77), .B1(new_n230_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT77), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n222_), .A2(new_n229_), .A3(new_n236_), .A4(new_n233_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n230_), .A2(KEYINPUT76), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n222_), .A2(new_n229_), .A3(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n234_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT80), .B(G176gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G169gat), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n245_), .A2(new_n246_), .B1(G169gat), .B2(G176gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G183gat), .A2(G190gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT23), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n250_), .B(new_n251_), .C1(G183gat), .C2(G190gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT25), .B(G183gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT78), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G183gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n257_), .B2(KEYINPUT25), .ZN(new_n258_));
  INV_X1    g057(.A(G190gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT26), .B1(new_n259_), .B2(KEYINPUT79), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT26), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(G190gat), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n258_), .B(new_n260_), .C1(KEYINPUT79), .C2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n256_), .A2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n250_), .A2(new_n251_), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G176gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(KEYINPUT24), .A3(new_n269_), .ZN(new_n270_));
  OR3_X1    g069(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n265_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n253_), .B1(new_n264_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT81), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT81), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n253_), .B(new_n275_), .C1(new_n264_), .C2(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278_));
  INV_X1    g077(.A(G43gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n277_), .B(new_n280_), .Z(new_n281_));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(new_n206_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT30), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT82), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n284_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G113gat), .B(G120gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n290_), .B(new_n291_), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT31), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n288_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT82), .B1(new_n295_), .B2(new_n285_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n289_), .A3(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT85), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT2), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT2), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(G141gat), .A3(G148gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n308_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT84), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n303_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n313_), .B(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(KEYINPUT83), .B(KEYINPUT3), .Z(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n310_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n317_), .A2(new_n319_), .A3(KEYINPUT85), .A4(new_n308_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n302_), .B1(new_n315_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n301_), .A2(KEYINPUT1), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(new_n299_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n301_), .A2(KEYINPUT1), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(new_n304_), .A3(new_n311_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n322_), .A2(new_n323_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT86), .B1(new_n321_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n331_), .A3(new_n292_), .ZN(new_n332_));
  OR3_X1    g131(.A1(new_n321_), .A2(new_n292_), .A3(new_n330_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT4), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n329_), .A2(new_n331_), .A3(new_n337_), .A4(new_n292_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n332_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G1gat), .B(G29gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(new_n340_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT27), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G8gat), .B(G36gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT18), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G64gat), .B(G92gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT89), .B(G204gat), .ZN(new_n355_));
  INV_X1    g154(.A(G197gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT21), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(G197gat), .B2(G204gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n355_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n367_));
  INV_X1    g166(.A(G204gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(G197gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n355_), .B2(G197gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n364_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n366_), .A2(new_n370_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n361_), .A2(new_n358_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n362_), .A2(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n355_), .A2(G197gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n369_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n365_), .A3(new_n373_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n363_), .B1(new_n379_), .B2(new_n365_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n360_), .A2(new_n361_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n265_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT26), .B(G190gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n254_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n253_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n376_), .B1(new_n383_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n375_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT19), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT93), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT93), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n390_), .A2(new_n395_), .A3(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n362_), .A2(new_n371_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n384_), .A2(new_n386_), .B1(new_n252_), .B2(new_n247_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n380_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT95), .ZN(new_n401_));
  INV_X1    g200(.A(new_n392_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT20), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n383_), .A2(new_n388_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT95), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n276_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n271_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n408_), .B(new_n270_), .C1(new_n256_), .C2(new_n263_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n275_), .B1(new_n409_), .B2(new_n253_), .ZN(new_n410_));
  OAI211_X1 g209(.A(KEYINPUT94), .B(new_n383_), .C1(new_n407_), .C2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT94), .B1(new_n277_), .B2(new_n383_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n401_), .B(new_n406_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n354_), .B1(new_n397_), .B2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n395_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n416_));
  AOI211_X1 g215(.A(KEYINPUT93), .B(new_n402_), .C1(new_n375_), .C2(new_n389_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n414_), .B(new_n354_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n350_), .B1(new_n415_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(KEYINPUT100), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT100), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n397_), .A2(new_n422_), .A3(new_n354_), .A4(new_n414_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n354_), .ZN(new_n424_));
  XOR2_X1   g223(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n425_));
  OAI211_X1 g224(.A(KEYINPUT98), .B(new_n425_), .C1(new_n383_), .C2(new_n388_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT98), .B1(new_n400_), .B2(new_n425_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n383_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT94), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n411_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n402_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n390_), .A2(new_n392_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n424_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n421_), .A2(new_n423_), .A3(KEYINPUT27), .A4(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n349_), .A2(new_n420_), .A3(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G22gat), .B(G50gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n329_), .A2(new_n331_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT29), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT87), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n446_));
  AOI211_X1 g245(.A(new_n446_), .B(KEYINPUT29), .C1(new_n329_), .C2(new_n331_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n442_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n331_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n321_), .A2(KEYINPUT86), .A3(new_n330_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n444_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n446_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n443_), .A2(KEYINPUT87), .A3(new_n444_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n441_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT92), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G228gat), .A2(G233gat), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n457_), .B(new_n383_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n444_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n459_));
  OAI211_X1 g258(.A(G228gat), .B(G233gat), .C1(new_n459_), .C2(new_n374_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G78gat), .B(G106gat), .Z(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n462_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n458_), .A2(new_n460_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n448_), .A2(new_n454_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n456_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n455_), .A2(KEYINPUT92), .A3(new_n463_), .A4(new_n465_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n438_), .A2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n415_), .A2(new_n419_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n339_), .A2(KEYINPUT33), .A3(new_n340_), .A4(new_n345_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n346_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n334_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n345_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n332_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n473_), .A2(new_n474_), .A3(new_n476_), .A4(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n332_), .A2(KEYINPUT4), .A3(new_n333_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n338_), .A2(new_n336_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n340_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n478_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n346_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n354_), .A2(KEYINPUT32), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n414_), .B(new_n487_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT99), .ZN(new_n489_));
  INV_X1    g288(.A(new_n487_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(KEYINPUT99), .B(new_n490_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n486_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n481_), .A2(new_n494_), .B1(new_n470_), .B2(new_n469_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n298_), .B1(new_n472_), .B2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n420_), .A2(new_n437_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n471_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n298_), .A2(new_n486_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n496_), .A2(KEYINPUT101), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT101), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n503_), .B(new_n298_), .C1(new_n472_), .C2(new_n495_), .ZN(new_n504_));
  AOI211_X1 g303(.A(KEYINPUT102), .B(new_n244_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT102), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n496_), .A2(KEYINPUT101), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n500_), .A2(new_n501_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n506_), .B1(new_n509_), .B2(new_n243_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511_));
  INV_X1    g310(.A(G99gat), .ZN(new_n512_));
  INV_X1    g311(.A(G106gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n514_), .A2(new_n517_), .A3(new_n518_), .A4(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(G85gat), .ZN(new_n521_));
  INV_X1    g320(.A(G92gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G85gat), .A2(G92gat), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n520_), .A2(KEYINPUT8), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT8), .B1(new_n520_), .B2(new_n525_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n529_));
  OR2_X1    g328(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n513_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n523_), .A2(KEYINPUT9), .A3(new_n524_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(G85gat), .A3(G92gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n517_), .A2(new_n536_), .A3(new_n518_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n529_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n517_), .A2(new_n536_), .A3(new_n518_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n539_), .A2(KEYINPUT66), .A3(new_n532_), .A4(new_n533_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G57gat), .B(G64gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G71gat), .B(G78gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n545_));
  INV_X1    g344(.A(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n544_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n528_), .A2(new_n541_), .A3(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT12), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n528_), .A2(new_n541_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n549_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n555_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AOI211_X1 g357(.A(KEYINPUT12), .B(new_n549_), .C1(new_n528_), .C2(new_n541_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n554_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT67), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n553_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n556_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(new_n549_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n550_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n563_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n554_), .B(KEYINPUT67), .C1(new_n558_), .C2(new_n559_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n562_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G120gat), .B(G148gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(G176gat), .B(G204gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT69), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n569_), .A2(new_n574_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n569_), .A2(KEYINPUT69), .A3(new_n574_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n578_), .A2(KEYINPUT13), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT13), .B1(new_n578_), .B2(new_n579_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n505_), .A2(new_n510_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT73), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT74), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT35), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT72), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n564_), .A2(new_n219_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n595_), .A2(new_n596_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n225_), .A2(new_n556_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT71), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n225_), .A2(new_n556_), .A3(new_n604_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n602_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n600_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n598_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n600_), .A2(new_n601_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n610_), .A2(new_n603_), .A3(new_n597_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n590_), .B(new_n592_), .C1(new_n609_), .C2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n605_), .A2(new_n606_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n602_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n608_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n611_), .B1(new_n615_), .B2(new_n597_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n589_), .A3(new_n588_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n612_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT37), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n612_), .A2(new_n617_), .A3(KEYINPUT37), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n549_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(new_n212_), .ZN(new_n625_));
  XOR2_X1   g424(.A(G127gat), .B(G155gat), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT16), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT17), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n629_), .A2(new_n630_), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n625_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n625_), .A2(new_n631_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n622_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n583_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n349_), .A2(G1gat), .ZN(new_n640_));
  OR3_X1    g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n612_), .A2(new_n617_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n582_), .A2(new_n244_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n643_), .A2(new_n635_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n486_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G1gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n639_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n641_), .A2(new_n647_), .A3(new_n648_), .ZN(G1324gat));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n645_), .A2(new_n498_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n652_), .B2(G8gat), .ZN(new_n653_));
  INV_X1    g452(.A(G8gat), .ZN(new_n654_));
  AOI211_X1 g453(.A(KEYINPUT39), .B(new_n654_), .C1(new_n645_), .C2(new_n498_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n498_), .A2(new_n654_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n638_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n650_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  OAI221_X1 g458(.A(KEYINPUT40), .B1(new_n638_), .B2(new_n657_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1325gat));
  INV_X1    g460(.A(new_n298_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n206_), .B1(new_n645_), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n206_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n638_), .B2(new_n665_), .ZN(G1326gat));
  AOI21_X1  g465(.A(new_n207_), .B1(new_n645_), .B2(new_n499_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT42), .Z(new_n668_));
  NAND2_X1  g467(.A1(new_n499_), .A2(new_n207_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n638_), .B2(new_n669_), .ZN(G1327gat));
  NOR2_X1   g469(.A1(new_n618_), .A2(new_n635_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n583_), .A2(new_n671_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n672_), .A2(G29gat), .A3(new_n349_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n644_), .A2(new_n636_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n621_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT37), .B1(new_n612_), .B2(new_n617_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT43), .B(new_n678_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n509_), .B2(new_n622_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT44), .B(new_n675_), .C1(new_n679_), .C2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n481_), .A2(new_n494_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n471_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n497_), .A2(new_n470_), .A3(new_n469_), .A4(new_n349_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n662_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n508_), .B1(new_n686_), .B2(new_n503_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n504_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n622_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT43), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n509_), .A2(new_n680_), .A3(new_n622_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n674_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n682_), .B(new_n486_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(new_n695_), .A3(G29gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n694_), .B2(G29gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n673_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  OAI211_X1 g497(.A(new_n682_), .B(new_n498_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n497_), .A2(G36gat), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n583_), .A2(new_n701_), .A3(new_n671_), .A4(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n243_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n582_), .B1(new_n704_), .B2(KEYINPUT102), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n509_), .A2(new_n506_), .A3(new_n243_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n671_), .A4(new_n702_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT45), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n703_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n700_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n700_), .A2(new_n709_), .A3(KEYINPUT46), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1329gat));
  XNOR2_X1  g513(.A(KEYINPUT105), .B(G43gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n715_), .B1(new_n672_), .B2(new_n298_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n298_), .A2(new_n279_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n682_), .B(new_n717_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT47), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n716_), .A2(new_n721_), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1330gat));
  INV_X1    g522(.A(G50gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n672_), .B2(new_n471_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n471_), .A2(new_n724_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n682_), .B(new_n726_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1331gat));
  INV_X1    g527(.A(new_n582_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n729_), .A2(new_n636_), .A3(new_n243_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n643_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n349_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n729_), .A2(new_n243_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n509_), .A2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(new_n637_), .ZN(new_n736_));
  INV_X1    g535(.A(G57gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n737_), .A3(new_n486_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n733_), .A2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n736_), .A2(new_n740_), .A3(new_n498_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n731_), .A2(new_n498_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G64gat), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT48), .B(new_n740_), .C1(new_n731_), .C2(new_n498_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT106), .ZN(G1333gat));
  INV_X1    g546(.A(G71gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n731_), .B2(new_n662_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT49), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n736_), .A2(new_n748_), .A3(new_n662_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n731_), .B2(new_n499_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT50), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n736_), .A2(new_n753_), .A3(new_n499_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1335gat));
  NAND3_X1  g556(.A1(new_n735_), .A2(new_n486_), .A3(new_n671_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n521_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(new_n521_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n690_), .A2(new_n691_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n734_), .A2(new_n636_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT108), .Z(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n486_), .A2(G85gat), .ZN(new_n766_));
  OAI22_X1  g565(.A1(new_n760_), .A2(new_n761_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(G1336gat));
  AND2_X1   g568(.A1(new_n735_), .A2(new_n671_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G92gat), .B1(new_n770_), .B2(new_n498_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n765_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n497_), .A2(new_n522_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT110), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n772_), .B2(new_n774_), .ZN(G1337gat));
  OAI21_X1  g574(.A(G99gat), .B1(new_n765_), .B2(new_n298_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n770_), .A2(new_n530_), .A3(new_n531_), .A4(new_n662_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n770_), .A2(new_n513_), .A3(new_n499_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n764_), .B(new_n499_), .C1(new_n681_), .C2(new_n679_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(new_n782_), .A3(G106gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G106gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT53), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(new_n780_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790_));
  NOR4_X1   g589(.A1(new_n498_), .A2(new_n499_), .A3(new_n298_), .A4(new_n349_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n560_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n550_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n563_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n795_), .B2(new_n563_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n562_), .A2(new_n793_), .A3(new_n568_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n574_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n574_), .A2(KEYINPUT56), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n800_), .B(new_n794_), .C1(new_n798_), .C2(new_n797_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(KEYINPUT114), .A3(new_n805_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n804_), .A2(new_n808_), .A3(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n202_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n223_), .A2(new_n228_), .A3(new_n203_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n234_), .A3(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n238_), .A2(new_n814_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n815_), .A2(new_n575_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT58), .B1(new_n811_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n792_), .B1(new_n817_), .B2(new_n678_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n575_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n807_), .A2(new_n806_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n810_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT115), .B(new_n622_), .C1(new_n821_), .C2(KEYINPUT58), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(KEYINPUT58), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n806_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n574_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n243_), .B(new_n575_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n815_), .A2(new_n579_), .A3(new_n578_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT57), .B1(new_n829_), .B2(new_n618_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  AOI211_X1 g630(.A(new_n831_), .B(new_n642_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n635_), .B1(new_n824_), .B2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n243_), .A2(new_n636_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT111), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n729_), .A2(new_n836_), .A3(new_n678_), .ZN(new_n837_));
  XOR2_X1   g636(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n729_), .A2(new_n836_), .A3(new_n678_), .A4(new_n838_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n791_), .B1(new_n834_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT59), .B(new_n791_), .C1(new_n834_), .C2(new_n842_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n845_), .A2(KEYINPUT116), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT116), .B1(new_n845_), .B2(new_n846_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n243_), .A2(G113gat), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n843_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n243_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n790_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n852_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n845_), .A2(new_n846_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n845_), .A2(KEYINPUT116), .A3(new_n846_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT117), .B(new_n854_), .C1(new_n859_), .C2(new_n849_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n853_), .A2(new_n860_), .ZN(G1340gat));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n729_), .B2(KEYINPUT60), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n851_), .B(new_n863_), .C1(KEYINPUT60), .C2(new_n862_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n729_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n862_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n851_), .B2(new_n635_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n859_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT119), .B(G127gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n635_), .A2(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT120), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n869_), .B1(new_n870_), .B2(new_n873_), .ZN(G1342gat));
  INV_X1    g673(.A(G134gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n843_), .B2(new_n618_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT121), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n678_), .A2(new_n875_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n870_), .B2(new_n878_), .ZN(G1343gat));
  OR2_X1    g678(.A1(new_n834_), .A2(new_n842_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n662_), .A2(new_n471_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n498_), .A2(new_n349_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n244_), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n729_), .ZN(new_n886_));
  XOR2_X1   g685(.A(KEYINPUT122), .B(G148gat), .Z(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1345gat));
  OR3_X1    g687(.A1(new_n883_), .A2(KEYINPUT123), .A3(new_n636_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT123), .B1(new_n883_), .B2(new_n636_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n883_), .B2(new_n678_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n618_), .A2(G162gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n883_), .B2(new_n896_), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n499_), .A2(new_n497_), .A3(new_n298_), .A4(new_n486_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n880_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n243_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n898_), .B1(new_n902_), .B2(new_n266_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n246_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(new_n904_), .A3(new_n905_), .ZN(G1348gat));
  NAND2_X1  g705(.A1(new_n900_), .A2(new_n582_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT125), .B1(new_n907_), .B2(new_n267_), .ZN(new_n908_));
  OR3_X1    g707(.A1(new_n907_), .A2(KEYINPUT125), .A3(new_n267_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n245_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n907_), .A2(KEYINPUT124), .A3(new_n245_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n908_), .A2(new_n909_), .B1(new_n912_), .B2(new_n913_), .ZN(G1349gat));
  NAND2_X1  g713(.A1(new_n900_), .A2(new_n635_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n254_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n257_), .B2(new_n915_), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n900_), .A2(new_n642_), .A3(new_n385_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n900_), .A2(new_n622_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n919_), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(KEYINPUT126), .B1(new_n919_), .B2(G190gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n918_), .B1(new_n920_), .B2(new_n921_), .ZN(G1351gat));
  NAND4_X1  g721(.A1(new_n880_), .A2(new_n349_), .A3(new_n498_), .A4(new_n881_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n244_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n356_), .ZN(G1352gat));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n729_), .ZN(new_n926_));
  MUX2_X1   g725(.A(G204gat), .B(new_n355_), .S(new_n926_), .Z(G1353gat));
  NAND2_X1  g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n635_), .A2(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(KEYINPUT127), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n923_), .A2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1354gat));
  OAI21_X1  g732(.A(G218gat), .B1(new_n923_), .B2(new_n678_), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n618_), .A2(G218gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n923_), .B2(new_n935_), .ZN(G1355gat));
endmodule


