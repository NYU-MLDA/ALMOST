//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n203_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT22), .B1(new_n211_), .B2(KEYINPUT82), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT82), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT22), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT83), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n217_), .A2(new_n218_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n210_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n205_), .A2(KEYINPUT81), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT81), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n204_), .B2(KEYINPUT23), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n207_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n202_), .A2(KEYINPUT24), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  MUX2_X1   g026(.A(new_n226_), .B(KEYINPUT24), .S(new_n227_), .Z(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT26), .B(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(G183gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT25), .B1(new_n230_), .B2(KEYINPUT80), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(KEYINPUT25), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n229_), .B(new_n231_), .C1(new_n232_), .C2(KEYINPUT80), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n225_), .A2(new_n228_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT84), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n221_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n221_), .B2(new_n234_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G99gat), .ZN(new_n239_));
  INV_X1    g038(.A(G43gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n238_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  INV_X1    g042(.A(G15gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT30), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n242_), .B(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n247_), .A2(KEYINPUT85), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(KEYINPUT85), .ZN(new_n249_));
  XOR2_X1   g048(.A(G127gat), .B(G134gat), .Z(new_n250_));
  XOR2_X1   g049(.A(G113gat), .B(G120gat), .Z(new_n251_));
  XOR2_X1   g050(.A(new_n250_), .B(new_n251_), .Z(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT31), .ZN(new_n253_));
  OR3_X1    g052(.A1(new_n248_), .A2(new_n249_), .A3(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n247_), .A2(KEYINPUT85), .A3(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G1gat), .B(G29gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT103), .B(G85gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G57gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  NAND2_X1  g061(.A1(G225gat), .A2(G233gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G141gat), .A2(G148gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT86), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(KEYINPUT1), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G155gat), .B(G162gat), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n268_), .B(new_n271_), .C1(KEYINPUT1), .C2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(KEYINPUT89), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT2), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n266_), .A2(new_n275_), .A3(new_n267_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n264_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT2), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n269_), .A2(KEYINPUT87), .A3(KEYINPUT3), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT3), .B1(new_n269_), .B2(KEYINPUT87), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n276_), .B(new_n278_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n274_), .B1(new_n282_), .B2(KEYINPUT88), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT88), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n269_), .A2(KEYINPUT87), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n287_), .A2(new_n279_), .B1(KEYINPUT2), .B2(new_n277_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n284_), .B1(new_n288_), .B2(new_n276_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n273_), .B1(new_n283_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n252_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n252_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n292_), .B(new_n273_), .C1(new_n283_), .C2(new_n289_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(KEYINPUT4), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n291_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n294_), .A2(KEYINPUT102), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT102), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n291_), .A2(new_n293_), .A3(new_n298_), .A4(KEYINPUT4), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n263_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n291_), .A2(new_n293_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n263_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n262_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n294_), .A2(KEYINPUT102), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n295_), .A2(new_n296_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n299_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n303_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n262_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n304_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n305_), .A2(new_n312_), .A3(KEYINPUT106), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT106), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n314_), .B(new_n262_), .C1(new_n300_), .C2(new_n304_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n257_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G197gat), .A2(G204gat), .ZN(new_n319_));
  INV_X1    g118(.A(G204gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT90), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT90), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G204gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n319_), .B1(new_n324_), .B2(G197gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT94), .ZN(new_n326_));
  XOR2_X1   g125(.A(G211gat), .B(G218gat), .Z(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(KEYINPUT21), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT92), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(new_n325_), .B2(KEYINPUT21), .ZN(new_n330_));
  INV_X1    g129(.A(new_n319_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT90), .B(G204gat), .ZN(new_n332_));
  INV_X1    g131(.A(G197gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT21), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT92), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(G197gat), .B2(G204gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n324_), .B2(G197gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT91), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(KEYINPUT91), .B(new_n338_), .C1(new_n324_), .C2(G197gat), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n327_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT93), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n337_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(new_n337_), .B2(new_n343_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n328_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n229_), .ZN(new_n348_));
  XOR2_X1   g147(.A(KEYINPUT25), .B(G183gat), .Z(new_n349_));
  OAI211_X1 g148(.A(new_n228_), .B(new_n208_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n225_), .A2(new_n209_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G169gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n203_), .B1(new_n352_), .B2(new_n216_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n351_), .A2(KEYINPUT98), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT98), .B1(new_n351_), .B2(new_n353_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n350_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n347_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT20), .ZN(new_n358_));
  INV_X1    g157(.A(new_n238_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n347_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n357_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT99), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n358_), .B1(new_n347_), .B2(new_n356_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n337_), .A2(new_n343_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT93), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n337_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n238_), .A3(new_n328_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n365_), .B1(new_n372_), .B2(new_n362_), .ZN(new_n373_));
  AOI211_X1 g172(.A(KEYINPUT99), .B(new_n363_), .C1(new_n366_), .C2(new_n371_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n364_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G8gat), .B(G36gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n380_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n382_), .B(new_n364_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(KEYINPUT101), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT101), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n375_), .A2(new_n386_), .A3(new_n380_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT96), .ZN(new_n389_));
  INV_X1    g188(.A(G228gat), .ZN(new_n390_));
  INV_X1    g189(.A(G233gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT95), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n347_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n370_), .A2(KEYINPUT95), .A3(new_n328_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n290_), .A2(KEYINPUT29), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n389_), .B(new_n392_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n392_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT96), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n397_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(new_n400_), .A3(new_n347_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  OR3_X1    g204(.A1(new_n290_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT28), .B1(new_n290_), .B2(KEYINPUT29), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G22gat), .B(G50gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n406_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G78gat), .B(G106gat), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(KEYINPUT97), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n405_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n402_), .A2(new_n417_), .A3(new_n404_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n351_), .A2(new_n353_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n394_), .A2(new_n395_), .A3(new_n350_), .A4(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n363_), .B1(new_n424_), .B2(new_n360_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n372_), .A2(new_n362_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n380_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n383_), .A2(KEYINPUT27), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n388_), .A2(new_n422_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT108), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n388_), .A2(new_n422_), .A3(KEYINPUT108), .A4(new_n428_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n318_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n384_), .A2(new_n387_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n310_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT33), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n302_), .A2(KEYINPUT104), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT104), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n263_), .B1(new_n301_), .B2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n262_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n297_), .A2(new_n263_), .A3(new_n299_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n437_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n436_), .B1(new_n443_), .B2(new_n435_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n382_), .A2(KEYINPUT32), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT105), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(KEYINPUT105), .B(new_n447_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n375_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n450_), .A2(new_n451_), .B1(new_n452_), .B2(new_n446_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n434_), .A2(new_n445_), .B1(new_n453_), .B2(new_n316_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT107), .B1(new_n454_), .B2(new_n421_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT107), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n451_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(new_n446_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n316_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n444_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n456_), .B(new_n422_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n388_), .A2(new_n428_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n422_), .A2(new_n316_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n455_), .A2(new_n461_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n433_), .B1(new_n465_), .B2(new_n256_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT79), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT71), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n468_), .A2(KEYINPUT71), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(KEYINPUT71), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n470_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477_));
  INV_X1    g276(.A(G1gat), .ZN(new_n478_));
  INV_X1    g277(.A(G8gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G8gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n476_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT15), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n476_), .B(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n484_), .B1(new_n486_), .B2(new_n483_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G229gat), .A2(G233gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n467_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n476_), .B(new_n483_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT78), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(new_n467_), .A3(new_n488_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G113gat), .B(G141gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G169gat), .B(G197gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  OR2_X1    g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n497_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G230gat), .A2(G233gat), .ZN(new_n502_));
  AND2_X1   g301(.A1(G71gat), .A2(G78gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(G71gat), .A2(G78gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(KEYINPUT11), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n506_), .B2(KEYINPUT11), .ZN(new_n509_));
  INV_X1    g308(.A(G64gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(G57gat), .ZN(new_n511_));
  INV_X1    g310(.A(G57gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G64gat), .ZN(new_n513_));
  AND4_X1   g312(.A1(new_n508_), .A2(new_n511_), .A3(new_n513_), .A4(KEYINPUT11), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n507_), .B1(new_n509_), .B2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n511_), .A2(new_n513_), .A3(KEYINPUT11), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT68), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n511_), .A2(new_n513_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT11), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n511_), .A2(new_n513_), .A3(new_n508_), .A4(KEYINPUT11), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n517_), .A2(new_n520_), .A3(new_n505_), .A4(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(G85gat), .A2(G92gat), .ZN(new_n524_));
  AND2_X1   g323(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n531_));
  INV_X1    g330(.A(G99gat), .ZN(new_n532_));
  INV_X1    g331(.A(G106gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n527_), .B1(new_n530_), .B2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OAI221_X1 g338(.A(new_n527_), .B1(KEYINPUT67), .B2(KEYINPUT8), .C1(new_n530_), .C2(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n528_), .B(KEYINPUT6), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT10), .B(G99gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT64), .B(G106gat), .Z(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT66), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT9), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(G92gat), .ZN(new_n548_));
  INV_X1    g347(.A(G85gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT65), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT65), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(G85gat), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n524_), .A2(new_n526_), .A3(new_n547_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n546_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(G92gat), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(KEYINPUT9), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n551_), .A2(G85gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n549_), .A2(KEYINPUT65), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n526_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(KEYINPUT9), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(KEYINPUT66), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n545_), .B1(new_n555_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n523_), .B1(new_n541_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n543_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT64), .B(G106gat), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n530_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n553_), .A2(new_n554_), .A3(new_n546_), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT66), .B1(new_n560_), .B2(new_n563_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n515_), .A2(new_n522_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n539_), .A4(new_n540_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n502_), .B1(new_n566_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n566_), .A2(KEYINPUT12), .A3(new_n574_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n523_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n575_), .B1(new_n580_), .B2(new_n502_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n587_), .A2(KEYINPUT69), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n581_), .A2(new_n586_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT13), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(KEYINPUT13), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n573_), .B(new_n483_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT75), .ZN(new_n598_));
  XOR2_X1   g397(.A(G127gat), .B(G155gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT17), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n597_), .B1(new_n598_), .B2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n603_), .A2(KEYINPUT17), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n605_), .B2(KEYINPUT74), .ZN(new_n608_));
  INV_X1    g407(.A(new_n603_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT75), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n606_), .B(new_n608_), .C1(new_n597_), .C2(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT76), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(KEYINPUT76), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT77), .Z(new_n616_));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n486_), .A2(new_n577_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT35), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n577_), .A2(new_n476_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n618_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n622_), .A2(new_n623_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n627_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(KEYINPUT72), .A3(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G190gat), .B(G218gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n617_), .B1(new_n630_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n628_), .A2(new_n633_), .A3(new_n629_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n617_), .A3(new_n634_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n637_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n635_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT37), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n616_), .A2(new_n645_), .ZN(new_n646_));
  NOR4_X1   g445(.A1(new_n466_), .A2(new_n501_), .A3(new_n594_), .A4(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n478_), .A3(new_n316_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT38), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n593_), .A2(new_n615_), .A3(new_n500_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT109), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n466_), .B2(new_n639_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n422_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n653_));
  AOI22_X1  g452(.A1(new_n653_), .A2(KEYINPUT107), .B1(new_n462_), .B2(new_n463_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n257_), .B1(new_n654_), .B2(new_n461_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT109), .B(new_n643_), .C1(new_n655_), .C2(new_n433_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n650_), .B1(new_n652_), .B2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n657_), .A2(new_n316_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n649_), .B1(new_n478_), .B2(new_n658_), .ZN(G1324gat));
  INV_X1    g458(.A(new_n462_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n647_), .A2(new_n479_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n657_), .A2(new_n660_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(G8gat), .ZN(new_n664_));
  AOI211_X1 g463(.A(KEYINPUT39), .B(new_n479_), .C1(new_n657_), .C2(new_n660_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT40), .B(new_n661_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1325gat));
  NAND3_X1  g469(.A1(new_n647_), .A2(new_n244_), .A3(new_n257_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n657_), .A2(new_n257_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n672_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT41), .B1(new_n672_), .B2(G15gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n673_), .B2(new_n674_), .ZN(G1326gat));
  INV_X1    g474(.A(G22gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n421_), .A2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT110), .Z(new_n678_));
  NAND2_X1  g477(.A1(new_n647_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n657_), .A2(new_n421_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(G22gat), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT42), .B(new_n676_), .C1(new_n657_), .C2(new_n421_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n682_), .B2(new_n683_), .ZN(G1327gat));
  INV_X1    g483(.A(new_n466_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n594_), .A2(new_n616_), .A3(new_n643_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n685_), .A2(KEYINPUT111), .A3(new_n500_), .A4(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n500_), .B(new_n686_), .C1(new_n655_), .C2(new_n433_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT111), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n316_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n466_), .B2(new_n645_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  INV_X1    g493(.A(new_n645_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n694_), .B(new_n695_), .C1(new_n655_), .C2(new_n433_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n616_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n500_), .A3(new_n593_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n702_), .B(new_n699_), .C1(new_n693_), .C2(new_n696_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n316_), .A2(G29gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n692_), .B1(new_n704_), .B2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n704_), .B2(new_n660_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n687_), .A2(new_n690_), .A3(new_n708_), .A4(new_n660_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n710_), .B(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n707_), .B1(new_n709_), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n710_), .B(new_n711_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n701_), .A2(new_n703_), .A3(new_n462_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n715_), .B(KEYINPUT46), .C1(new_n716_), .C2(new_n708_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n717_), .ZN(G1329gat));
  AOI21_X1  g517(.A(G43gat), .B1(new_n691_), .B2(new_n257_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n256_), .A2(new_n240_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n704_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NOR4_X1   g522(.A1(new_n701_), .A2(new_n703_), .A3(new_n240_), .A4(new_n256_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT47), .B1(new_n724_), .B2(new_n719_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1330gat));
  INV_X1    g525(.A(G50gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n691_), .A2(new_n727_), .A3(new_n421_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n704_), .A2(new_n729_), .A3(new_n421_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G50gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n704_), .B2(new_n421_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1331gat));
  NOR4_X1   g532(.A1(new_n466_), .A2(new_n500_), .A3(new_n593_), .A4(new_n646_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n512_), .A3(new_n316_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n652_), .A2(new_n656_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n593_), .A2(new_n500_), .ZN(new_n737_));
  AND4_X1   g536(.A1(new_n316_), .A2(new_n736_), .A3(new_n616_), .A4(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n738_), .B2(new_n512_), .ZN(G1332gat));
  NAND3_X1  g538(.A1(new_n734_), .A2(new_n510_), .A3(new_n660_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n736_), .A2(new_n660_), .A3(new_n616_), .A4(new_n737_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G64gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n734_), .A2(new_n746_), .A3(new_n257_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n736_), .A2(new_n257_), .A3(new_n616_), .A4(new_n737_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(G71gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G71gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n734_), .A2(new_n753_), .A3(new_n421_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n736_), .A2(new_n421_), .A3(new_n616_), .A4(new_n737_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(G78gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G78gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n616_), .A2(new_n643_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n685_), .A2(KEYINPUT114), .A3(new_n760_), .A4(new_n737_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n760_), .B(new_n737_), .C1(new_n655_), .C2(new_n433_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n316_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n697_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n698_), .A2(new_n737_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n317_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(G1336gat));
  NAND3_X1  g570(.A1(new_n765_), .A2(new_n556_), .A3(new_n660_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n767_), .A2(new_n462_), .A3(new_n768_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(new_n556_), .ZN(G1337gat));
  NAND3_X1  g573(.A1(new_n765_), .A2(new_n257_), .A3(new_n567_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n767_), .A2(new_n256_), .A3(new_n768_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n532_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g577(.A(new_n768_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n697_), .A2(new_n421_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G106gat), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n422_), .A2(new_n544_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n765_), .A2(KEYINPUT115), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT115), .B1(new_n765_), .B2(new_n786_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT53), .B1(new_n785_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n789_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n787_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n784_), .A4(new_n783_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(new_n795_), .ZN(G1339gat));
  NAND4_X1  g595(.A1(new_n616_), .A2(new_n593_), .A3(new_n645_), .A4(new_n501_), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT54), .Z(new_n798_));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799_));
  INV_X1    g598(.A(new_n502_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n576_), .A2(new_n800_), .A3(new_n579_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n576_), .A2(KEYINPUT116), .A3(new_n800_), .A4(new_n579_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n580_), .B2(new_n502_), .ZN(new_n807_));
  AOI211_X1 g606(.A(KEYINPUT55), .B(new_n800_), .C1(new_n576_), .C2(new_n579_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n805_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT117), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n580_), .A2(new_n502_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT55), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n580_), .A2(new_n806_), .A3(new_n502_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n805_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n586_), .B1(new_n810_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n799_), .B1(new_n817_), .B2(KEYINPUT56), .ZN(new_n818_));
  AOI221_X4 g617(.A(KEYINPUT117), .B1(new_n803_), .B2(new_n804_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n815_), .B1(new_n814_), .B2(new_n805_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n585_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(KEYINPUT119), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n817_), .A2(KEYINPUT56), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n818_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n488_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n491_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(new_n497_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n487_), .A2(new_n826_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n494_), .A2(new_n497_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n830_), .A2(new_n587_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n825_), .A2(KEYINPUT58), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT120), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n825_), .A2(new_n831_), .A3(new_n834_), .A4(KEYINPUT58), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT58), .B1(new_n825_), .B2(new_n831_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n645_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT121), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n836_), .A2(new_n841_), .A3(new_n838_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n498_), .A2(new_n499_), .B1(new_n581_), .B2(new_n586_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n821_), .A2(new_n822_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n817_), .A2(KEYINPUT56), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n590_), .A2(new_n830_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n639_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n840_), .A2(new_n842_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n615_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n798_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n431_), .A2(new_n432_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n316_), .A3(new_n257_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT59), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(KEYINPUT59), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n616_), .B1(new_n839_), .B2(new_n850_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n797_), .B(KEYINPUT54), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n857_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n856_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G113gat), .B1(new_n864_), .B2(new_n501_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n853_), .A2(new_n855_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n501_), .A2(G113gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n865_), .B1(new_n867_), .B2(new_n868_), .ZN(G1340gat));
  OAI21_X1  g668(.A(KEYINPUT123), .B1(new_n864_), .B2(new_n593_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n856_), .A2(new_n863_), .A3(new_n871_), .A4(new_n594_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(G120gat), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(G120gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n593_), .B2(KEYINPUT60), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n866_), .B(new_n875_), .C1(KEYINPUT60), .C2(new_n874_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(G1341gat));
  OAI21_X1  g676(.A(G127gat), .B1(new_n864_), .B2(new_n852_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n698_), .A2(G127gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n867_), .B2(new_n879_), .ZN(G1342gat));
  INV_X1    g679(.A(G134gat), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n864_), .A2(new_n881_), .A3(new_n645_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n867_), .B2(new_n643_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT124), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n885_), .B(new_n881_), .C1(new_n867_), .C2(new_n643_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n882_), .B1(new_n884_), .B2(new_n886_), .ZN(G1343gat));
  INV_X1    g686(.A(new_n853_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n257_), .A2(new_n422_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n888_), .A2(new_n316_), .A3(new_n462_), .A4(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n501_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT125), .B(G141gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1344gat));
  OR3_X1    g692(.A1(new_n890_), .A2(G148gat), .A3(new_n593_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G148gat), .B1(new_n890_), .B2(new_n593_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1345gat));
  NOR2_X1   g695(.A1(new_n890_), .A2(new_n698_), .ZN(new_n897_));
  XOR2_X1   g696(.A(KEYINPUT61), .B(G155gat), .Z(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1346gat));
  OAI21_X1  g698(.A(G162gat), .B1(new_n890_), .B2(new_n645_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n643_), .A2(G162gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n890_), .B2(new_n901_), .ZN(G1347gat));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n860_), .A2(new_n862_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n462_), .A2(new_n316_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n257_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n421_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n501_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n903_), .B1(new_n909_), .B2(new_n211_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n352_), .ZN(new_n911_));
  OAI211_X1 g710(.A(KEYINPUT62), .B(G169gat), .C1(new_n908_), .C2(new_n501_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(G1348gat));
  INV_X1    g712(.A(new_n908_), .ZN(new_n914_));
  AOI21_X1  g713(.A(G176gat), .B1(new_n914_), .B2(new_n594_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n853_), .B2(new_n421_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n849_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n848_), .B(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(KEYINPUT121), .B2(new_n839_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n615_), .B1(new_n920_), .B2(new_n842_), .ZN(new_n921_));
  OAI211_X1 g720(.A(KEYINPUT126), .B(new_n422_), .C1(new_n921_), .C2(new_n798_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n917_), .A2(new_n922_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n906_), .A2(new_n216_), .A3(new_n593_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n915_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  NAND4_X1  g724(.A1(new_n904_), .A2(new_n349_), .A3(new_n615_), .A4(new_n907_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n905_), .A2(new_n257_), .A3(new_n616_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n927_), .B1(new_n917_), .B2(new_n922_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n928_), .B2(G183gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT127), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n931_), .B(new_n926_), .C1(new_n928_), .C2(G183gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1350gat));
  OAI21_X1  g732(.A(G190gat), .B1(new_n908_), .B2(new_n645_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n639_), .A2(new_n229_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n908_), .B2(new_n935_), .ZN(G1351gat));
  NAND3_X1  g735(.A1(new_n888_), .A2(new_n889_), .A3(new_n905_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n501_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n333_), .ZN(G1352gat));
  NOR3_X1   g738(.A1(new_n937_), .A2(new_n332_), .A3(new_n593_), .ZN(new_n940_));
  OR2_X1    g739(.A1(new_n937_), .A2(new_n593_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n320_), .B2(new_n941_), .ZN(G1353gat));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  AND2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  NOR4_X1   g743(.A1(new_n937_), .A2(new_n852_), .A3(new_n943_), .A4(new_n944_), .ZN(new_n945_));
  OR2_X1    g744(.A1(new_n937_), .A2(new_n852_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(new_n943_), .ZN(G1354gat));
  OAI21_X1  g746(.A(G218gat), .B1(new_n937_), .B2(new_n645_), .ZN(new_n948_));
  OR2_X1    g747(.A1(new_n643_), .A2(G218gat), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n937_), .B2(new_n949_), .ZN(G1355gat));
endmodule


