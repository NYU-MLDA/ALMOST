//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n963_, new_n964_, new_n965_,
    new_n967_, new_n968_, new_n969_, new_n971_, new_n972_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  AND2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT82), .B(G176gat), .Z(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT22), .B(G169gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  AND3_X1   g008(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(G183gat), .B2(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT93), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(G183gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT25), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n215_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(KEYINPUT25), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(G183gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT93), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n221_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT94), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228_));
  OR3_X1    g027(.A1(new_n206_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n225_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT95), .ZN(new_n232_));
  NOR4_X1   g031(.A1(new_n231_), .A2(new_n210_), .A3(new_n211_), .A4(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n228_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT95), .B1(new_n212_), .B2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n226_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n214_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G197gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G204gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT89), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(new_n240_), .A3(G204gat), .ZN(new_n244_));
  INV_X1    g043(.A(G204gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G197gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G218gat), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n248_), .A2(G211gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(G211gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n251_), .A3(KEYINPUT21), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT90), .ZN(new_n253_));
  INV_X1    g052(.A(new_n251_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT88), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G197gat), .B(G204gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT21), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n242_), .A2(new_n244_), .A3(new_n257_), .A4(new_n246_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n241_), .A2(new_n246_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(KEYINPUT88), .A3(KEYINPUT21), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n254_), .A2(new_n258_), .A3(new_n259_), .A4(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT90), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n247_), .A2(new_n251_), .A3(new_n263_), .A4(KEYINPUT21), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n253_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n205_), .B1(new_n239_), .B2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT80), .B(G190gat), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(KEYINPUT26), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n222_), .A2(new_n223_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT81), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT26), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(KEYINPUT26), .B2(G190gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT81), .ZN(new_n276_));
  INV_X1    g075(.A(new_n270_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n271_), .A2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n229_), .A2(new_n212_), .A3(new_n234_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n212_), .B1(G183gat), .B2(new_n268_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n279_), .A2(new_n280_), .B1(new_n209_), .B2(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n253_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT20), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n266_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n276_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n286_));
  NOR3_X1   g085(.A1(new_n269_), .A2(KEYINPUT81), .A3(new_n270_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n280_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n209_), .A2(new_n281_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT20), .B1(new_n290_), .B2(new_n265_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n238_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(new_n230_), .A3(new_n236_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n283_), .B1(new_n293_), .B2(new_n214_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n204_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT96), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n239_), .A2(new_n265_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT96), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(new_n204_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n285_), .B1(new_n296_), .B2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G8gat), .B(G36gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(G64gat), .B(G92gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n202_), .B1(new_n303_), .B2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n265_), .B1(new_n239_), .B2(KEYINPUT100), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT100), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n293_), .A2(new_n312_), .A3(new_n214_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n284_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT101), .B1(new_n316_), .B2(new_n204_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n298_), .A2(new_n205_), .A3(new_n299_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n284_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(new_n205_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n317_), .B1(new_n320_), .B2(KEYINPUT101), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n310_), .B(KEYINPUT103), .C1(new_n321_), .C2(new_n309_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT103), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n205_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n318_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT101), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT101), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(new_n319_), .B2(new_n205_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n309_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n285_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n301_), .B1(new_n300_), .B2(new_n204_), .ZN(new_n331_));
  AOI211_X1 g130(.A(KEYINPUT96), .B(new_n205_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n309_), .B(new_n330_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT27), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n323_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n322_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G141gat), .ZN(new_n342_));
  INV_X1    g141(.A(G148gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  OAI22_X1  g145(.A1(new_n344_), .A2(KEYINPUT3), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT86), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n348_), .A2(KEYINPUT86), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n347_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n345_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n341_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n353_), .A2(new_n354_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n344_), .ZN(new_n358_));
  OAI211_X1 g157(.A(KEYINPUT85), .B(new_n337_), .C1(new_n339_), .C2(KEYINPUT1), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n337_), .A2(KEYINPUT1), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n337_), .B1(new_n339_), .B2(KEYINPUT1), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n358_), .B1(new_n359_), .B2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n356_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n265_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n265_), .A2(KEYINPUT87), .B1(G228gat), .B2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n350_), .A2(new_n349_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n347_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n355_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n340_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n363_), .A2(new_n359_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n357_), .A3(new_n344_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT28), .B1(new_n377_), .B2(KEYINPUT29), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT28), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n365_), .A2(new_n379_), .A3(new_n366_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G22gat), .B(G50gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n384_), .B(KEYINPUT91), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n382_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n378_), .A2(new_n380_), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n383_), .A2(new_n388_), .B1(KEYINPUT92), .B2(new_n386_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n370_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n383_), .A2(new_n388_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n386_), .A2(KEYINPUT92), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n369_), .A3(new_n389_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT104), .B(KEYINPUT27), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n308_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n402_), .B2(new_n333_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405_));
  INV_X1    g204(.A(G43gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n290_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n282_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(G15gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT30), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT31), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n408_), .A2(new_n410_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT83), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n408_), .A2(new_n410_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n415_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n408_), .A2(new_n410_), .A3(new_n415_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(G127gat), .B(G134gat), .Z(new_n425_));
  XOR2_X1   g224(.A(G113gat), .B(G120gat), .Z(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n418_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(new_n418_), .B2(new_n424_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT102), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n428_), .B1(new_n356_), .B2(new_n364_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n374_), .A2(new_n376_), .A3(new_n427_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n433_), .A2(new_n434_), .A3(KEYINPUT4), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT98), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT98), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n433_), .A2(new_n434_), .A3(new_n441_), .A4(KEYINPUT4), .ZN(new_n442_));
  INV_X1    g241(.A(new_n433_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n438_), .B1(new_n446_), .B2(new_n437_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G1gat), .B(G29gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(G85gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT0), .B(G57gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n447_), .A2(new_n452_), .ZN(new_n453_));
  AOI211_X1 g252(.A(new_n451_), .B(new_n438_), .C1(new_n446_), .C2(new_n437_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n432_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n447_), .A2(new_n452_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n439_), .A2(KEYINPUT98), .B1(new_n443_), .B2(new_n444_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n436_), .B1(new_n457_), .B2(new_n442_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n451_), .B1(new_n458_), .B2(new_n438_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(new_n459_), .A3(KEYINPUT102), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n431_), .A2(new_n455_), .A3(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n336_), .A2(new_n398_), .A3(new_n404_), .A4(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT105), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n403_), .B1(new_n322_), .B2(new_n335_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n465_), .A2(KEYINPUT105), .A3(new_n398_), .A4(new_n461_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n455_), .A2(new_n397_), .A3(new_n460_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n326_), .A2(new_n328_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n308_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT103), .B1(new_n469_), .B2(new_n310_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n329_), .A2(new_n334_), .A3(new_n323_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n467_), .B(new_n404_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n451_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n473_), .B1(new_n446_), .B2(new_n437_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT99), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT99), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n473_), .B(new_n476_), .C1(new_n446_), .C2(new_n437_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n402_), .A3(new_n333_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n453_), .A2(KEYINPUT33), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n459_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n309_), .A2(KEYINPUT32), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n484_), .ZN(new_n486_));
  OAI22_X1  g285(.A1(new_n453_), .A2(new_n454_), .B1(new_n401_), .B2(new_n486_), .ZN(new_n487_));
  OAI22_X1  g286(.A1(new_n479_), .A2(new_n483_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n398_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n472_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n431_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n464_), .A2(new_n466_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G29gat), .B(G36gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G43gat), .B(G50gat), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT79), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502_));
  INV_X1    g301(.A(G1gat), .ZN(new_n503_));
  INV_X1    g302(.A(G8gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT14), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G1gat), .B(G8gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  XNOR2_X1  g307(.A(new_n501_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n501_), .A2(new_n508_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n499_), .B(KEYINPUT15), .ZN(new_n514_));
  INV_X1    g313(.A(new_n508_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n513_), .A2(new_n516_), .A3(new_n510_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G113gat), .B(G141gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(G169gat), .B(G197gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n518_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n492_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G230gat), .A2(G233gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(KEYINPUT64), .Z(new_n526_));
  OR3_X1    g325(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT6), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n527_), .B(new_n528_), .C1(new_n530_), .C2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G85gat), .B(G92gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT8), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT8), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n538_), .A3(new_n535_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT10), .ZN(new_n540_));
  INV_X1    g339(.A(G99gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(G106gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT65), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n542_), .A2(KEYINPUT65), .A3(new_n543_), .A4(new_n544_), .ZN(new_n548_));
  INV_X1    g347(.A(G85gat), .ZN(new_n549_));
  INV_X1    g348(.A(G92gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(KEYINPUT9), .ZN(new_n551_));
  OR2_X1    g350(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .A4(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n547_), .A2(new_n548_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n554_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n531_), .A2(KEYINPUT6), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n529_), .A2(G99gat), .A3(G106gat), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n557_), .A2(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n537_), .A2(new_n539_), .B1(new_n556_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(G64gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(G57gat), .ZN(new_n564_));
  INV_X1    g363(.A(G57gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(G64gat), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n564_), .A2(new_n566_), .A3(KEYINPUT67), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT67), .B1(new_n564_), .B2(new_n566_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT11), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT67), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n565_), .A2(G64gat), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n563_), .A2(G57gat), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT11), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n564_), .A2(new_n566_), .A3(KEYINPUT67), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(G78gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(G71gat), .ZN(new_n578_));
  INV_X1    g377(.A(G71gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(G78gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n569_), .A2(new_n576_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n573_), .A2(new_n575_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n581_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(KEYINPUT11), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n562_), .A2(new_n586_), .ZN(new_n587_));
  AOI211_X1 g386(.A(new_n574_), .B(new_n581_), .C1(new_n573_), .C2(new_n575_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n584_), .B1(new_n583_), .B2(KEYINPUT11), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n589_), .B2(new_n576_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n561_), .A2(new_n548_), .A3(new_n555_), .A4(new_n547_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n528_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n559_), .A2(new_n560_), .ZN(new_n595_));
  AOI211_X1 g394(.A(KEYINPUT8), .B(new_n534_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n538_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n591_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n590_), .A2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n526_), .B1(new_n587_), .B2(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT68), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT12), .B1(new_n590_), .B2(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n590_), .A2(new_n598_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT69), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n582_), .A2(new_n605_), .A3(new_n585_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n607_), .A2(KEYINPUT12), .A3(new_n608_), .A4(new_n598_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n526_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n604_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n600_), .A2(KEYINPUT68), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n601_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(G120gat), .B(G148gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT70), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n613_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n601_), .A2(new_n619_), .A3(new_n611_), .A4(new_n612_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n625_));
  NOR2_X1   g424(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(KEYINPUT72), .B2(KEYINPUT13), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT73), .ZN(new_n630_));
  INV_X1    g429(.A(new_n608_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(new_n606_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n508_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n632_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G127gat), .B(G155gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT16), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G183gat), .B(G211gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT17), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT78), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n635_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n634_), .A2(new_n586_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n634_), .A2(new_n586_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n639_), .B(KEYINPUT17), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n642_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(G232gat), .A2(G233gat), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT34), .Z(new_n649_));
  INV_X1    g448(.A(KEYINPUT35), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT75), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n514_), .A2(new_n598_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n649_), .A2(new_n650_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT74), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n499_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n598_), .B2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n654_), .B1(new_n655_), .B2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n652_), .A2(new_n653_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(G190gat), .B(G218gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(G134gat), .B(G162gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT36), .Z(new_n668_));
  AND3_X1   g467(.A1(new_n663_), .A2(new_n664_), .A3(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n667_), .A2(KEYINPUT36), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n669_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT37), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT76), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n663_), .A2(new_n664_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n670_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n663_), .A2(new_n664_), .A3(new_n668_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT76), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(KEYINPUT37), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n677_), .A2(new_n674_), .A3(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT77), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT77), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n677_), .A2(new_n684_), .A3(new_n674_), .A4(new_n678_), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n675_), .A2(new_n681_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AND4_X1   g486(.A1(new_n524_), .A2(new_n630_), .A3(new_n647_), .A4(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n455_), .A2(new_n460_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n503_), .A3(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n691_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n679_), .A2(KEYINPUT107), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n679_), .A2(KEYINPUT107), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n492_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n647_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n629_), .A2(new_n523_), .A3(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n689_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G1gat), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n692_), .A2(new_n693_), .A3(new_n704_), .ZN(G1324gat));
  INV_X1    g504(.A(new_n465_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n688_), .A2(new_n504_), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT39), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n701_), .A2(new_n706_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(G8gat), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT39), .B(new_n504_), .C1(new_n701_), .C2(new_n706_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT40), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(G1325gat));
  NAND3_X1  g513(.A1(new_n688_), .A2(new_n412_), .A3(new_n431_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT108), .Z(new_n716_));
  OAI21_X1  g515(.A(G15gat), .B1(new_n702_), .B2(new_n491_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT41), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n717_), .A2(KEYINPUT41), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(new_n718_), .A3(new_n719_), .ZN(G1326gat));
  INV_X1    g519(.A(G22gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n701_), .B2(new_n397_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT42), .Z(new_n723_));
  NAND3_X1  g522(.A1(new_n688_), .A2(new_n721_), .A3(new_n397_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1327gat));
  NAND2_X1  g524(.A1(new_n673_), .A2(new_n699_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n629_), .A2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n524_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G29gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n689_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n464_), .A2(new_n466_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n431_), .B1(new_n472_), .B2(new_n489_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n731_), .B(new_n686_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n492_), .B2(new_n687_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n627_), .A2(new_n628_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n522_), .A3(new_n699_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT44), .B1(new_n736_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n741_), .B(new_n738_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n689_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G29gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n743_), .B2(new_n689_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n730_), .B1(new_n746_), .B2(new_n747_), .ZN(G1328gat));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  INV_X1    g548(.A(G36gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n743_), .B2(new_n706_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n728_), .A2(new_n750_), .A3(new_n706_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT111), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n752_), .B(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n749_), .B1(new_n751_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n752_), .B(new_n754_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n740_), .A2(new_n742_), .A3(new_n465_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n758_), .B(KEYINPUT46), .C1(new_n750_), .C2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(G1329gat));
  AOI21_X1  g560(.A(G43gat), .B1(new_n728_), .B2(new_n431_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n491_), .A2(new_n406_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n743_), .B2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(KEYINPUT47), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n766_), .B(new_n762_), .C1(new_n743_), .C2(new_n763_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1330gat));
  NAND2_X1  g567(.A1(new_n397_), .A2(G50gat), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n740_), .A2(new_n742_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771_));
  AOI21_X1  g570(.A(G50gat), .B1(new_n728_), .B2(new_n397_), .ZN(new_n772_));
  OR3_X1    g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n771_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1331gat));
  NOR2_X1   g574(.A1(new_n492_), .A2(new_n522_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n686_), .A2(new_n737_), .A3(new_n699_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n778_), .A2(G57gat), .A3(new_n703_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n523_), .A2(new_n647_), .ZN(new_n780_));
  NOR4_X1   g579(.A1(new_n492_), .A2(new_n630_), .A3(new_n697_), .A4(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n565_), .B1(new_n781_), .B2(new_n689_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT113), .ZN(G1332gat));
  AOI21_X1  g583(.A(new_n563_), .B1(new_n781_), .B2(new_n706_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT48), .Z(new_n786_));
  INV_X1    g585(.A(new_n778_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n563_), .A3(new_n706_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1333gat));
  NAND3_X1  g588(.A1(new_n787_), .A2(new_n579_), .A3(new_n431_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n781_), .A2(new_n431_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G71gat), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT49), .B(new_n579_), .C1(new_n781_), .C2(new_n431_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT114), .ZN(G1334gat));
  AOI21_X1  g595(.A(new_n577_), .B1(new_n781_), .B2(new_n397_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n797_), .B(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n787_), .A2(new_n577_), .A3(new_n397_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1335gat));
  NOR4_X1   g600(.A1(new_n492_), .A2(new_n630_), .A3(new_n522_), .A4(new_n726_), .ZN(new_n802_));
  AOI21_X1  g601(.A(G85gat), .B1(new_n802_), .B2(new_n689_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT116), .ZN(new_n804_));
  INV_X1    g603(.A(new_n736_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n522_), .A2(new_n647_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n629_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n703_), .A2(new_n549_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n804_), .B1(new_n808_), .B2(new_n809_), .ZN(G1336gat));
  NAND3_X1  g609(.A1(new_n802_), .A2(new_n550_), .A3(new_n706_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n805_), .A2(new_n465_), .A3(new_n807_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n550_), .ZN(G1337gat));
  NAND4_X1  g612(.A1(new_n802_), .A2(new_n431_), .A3(new_n542_), .A4(new_n544_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n805_), .A2(new_n491_), .A3(new_n807_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n541_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g616(.A1(new_n802_), .A2(new_n543_), .A3(new_n397_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n736_), .A2(new_n397_), .A3(new_n629_), .A4(new_n806_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n543_), .B1(new_n820_), .B2(KEYINPUT52), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(KEYINPUT52), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n819_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n818_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT53), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n827_), .B(new_n818_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1339gat));
  NAND4_X1  g628(.A1(new_n687_), .A2(new_n523_), .A3(new_n737_), .A4(new_n647_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT54), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n613_), .A2(new_n618_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n522_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n604_), .A2(new_n610_), .A3(new_n609_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n610_), .B1(new_n604_), .B2(new_n609_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n604_), .A2(new_n609_), .A3(new_n837_), .A4(new_n610_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT118), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT12), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n562_), .B2(new_n586_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n587_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n598_), .A2(KEYINPUT12), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n845_), .A2(new_n631_), .A3(new_n606_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n526_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(KEYINPUT55), .A3(new_n611_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n839_), .ZN(new_n850_));
  AND4_X1   g649(.A1(KEYINPUT56), .A2(new_n841_), .A3(new_n618_), .A4(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n618_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n839_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(KEYINPUT118), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT56), .B1(new_n854_), .B2(new_n850_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n834_), .B1(new_n851_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n521_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n513_), .A2(new_n516_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT119), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n511_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(KEYINPUT119), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n858_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n512_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n623_), .A2(new_n857_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n857_), .B1(new_n623_), .B2(new_n866_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n673_), .B1(new_n856_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n832_), .A2(new_n866_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n841_), .A2(new_n618_), .A3(new_n850_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT56), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n854_), .A2(KEYINPUT56), .A3(new_n850_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n871_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n686_), .B1(new_n876_), .B2(KEYINPUT58), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n878_), .B(new_n871_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n879_));
  OAI22_X1  g678(.A1(KEYINPUT57), .A2(new_n870_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT121), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n876_), .A2(KEYINPUT58), .ZN(new_n882_));
  INV_X1    g681(.A(new_n879_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(new_n883_), .A3(new_n686_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n833_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n868_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n623_), .A2(new_n857_), .A3(new_n866_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n679_), .B1(new_n885_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n884_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n889_), .A2(new_n890_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n881_), .A2(new_n893_), .A3(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n831_), .B1(new_n896_), .B2(new_n647_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n706_), .A2(new_n703_), .A3(new_n397_), .A4(new_n491_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n699_), .B1(new_n880_), .B2(new_n894_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n831_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n899_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT59), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n900_), .A2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G113gat), .B1(new_n905_), .B2(new_n523_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n523_), .A2(G113gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n903_), .B2(new_n907_), .ZN(G1340gat));
  XNOR2_X1  g707(.A(KEYINPUT122), .B(G120gat), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n910_), .B1(new_n905_), .B2(new_n630_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n909_), .A2(KEYINPUT60), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n909_), .B1(new_n737_), .B2(KEYINPUT60), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n902_), .A2(new_n899_), .A3(new_n912_), .A4(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT123), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n911_), .A2(new_n915_), .ZN(G1341gat));
  OAI21_X1  g715(.A(G127gat), .B1(new_n905_), .B2(new_n699_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n699_), .A2(G127gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n903_), .B2(new_n918_), .ZN(G1342gat));
  OAI21_X1  g718(.A(G134gat), .B1(new_n905_), .B2(new_n687_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n696_), .A2(G134gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n903_), .B2(new_n921_), .ZN(G1343gat));
  AOI21_X1  g721(.A(new_n431_), .B1(new_n831_), .B2(new_n901_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n706_), .A2(new_n703_), .A3(new_n398_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n523_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT124), .B(G141gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1344gat));
  NOR2_X1   g727(.A1(new_n925_), .A2(new_n630_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n343_), .ZN(G1345gat));
  OR3_X1    g729(.A1(new_n925_), .A2(KEYINPUT125), .A3(new_n699_), .ZN(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT125), .B1(new_n925_), .B2(new_n699_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(KEYINPUT61), .B(G155gat), .ZN(new_n933_));
  AND3_X1   g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1346gat));
  OAI21_X1  g735(.A(G162gat), .B1(new_n925_), .B2(new_n687_), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n696_), .A2(G162gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n925_), .B2(new_n938_), .ZN(G1347gat));
  NAND2_X1  g738(.A1(new_n706_), .A2(new_n461_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n397_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n894_), .B1(new_n880_), .B2(KEYINPUT121), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n647_), .B1(new_n942_), .B2(new_n893_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n831_), .ZN(new_n944_));
  OAI211_X1 g743(.A(new_n522_), .B(new_n941_), .C1(new_n943_), .C2(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n945_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n897_), .A2(new_n208_), .A3(new_n522_), .A4(new_n941_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(KEYINPUT62), .B1(new_n945_), .B2(G169gat), .ZN(new_n949_));
  OAI21_X1  g748(.A(KEYINPUT126), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n945_), .A2(G169gat), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n953_), .A2(new_n954_), .A3(new_n947_), .A4(new_n946_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n950_), .A2(new_n955_), .ZN(G1348gat));
  AND2_X1   g755(.A1(new_n897_), .A2(new_n941_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n629_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n397_), .B1(new_n831_), .B2(new_n901_), .ZN(new_n959_));
  INV_X1    g758(.A(G176gat), .ZN(new_n960_));
  NOR3_X1   g759(.A1(new_n630_), .A2(new_n960_), .A3(new_n940_), .ZN(new_n961_));
  AOI22_X1  g760(.A1(new_n958_), .A2(new_n207_), .B1(new_n959_), .B2(new_n961_), .ZN(G1349gat));
  NOR2_X1   g761(.A1(new_n940_), .A2(new_n699_), .ZN(new_n963_));
  AOI21_X1  g762(.A(G183gat), .B1(new_n959_), .B2(new_n963_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n699_), .B1(new_n220_), .B2(new_n224_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n964_), .B1(new_n957_), .B2(new_n965_), .ZN(G1350gat));
  NAND2_X1  g765(.A1(new_n957_), .A2(new_n686_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n967_), .A2(G190gat), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n957_), .A2(new_n221_), .A3(new_n697_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1351gat));
  NAND3_X1  g769(.A1(new_n923_), .A2(new_n467_), .A3(new_n706_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n971_), .A2(new_n523_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(new_n240_), .ZN(G1352gat));
  NOR2_X1   g772(.A1(new_n971_), .A2(new_n630_), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n974_), .B1(new_n975_), .B2(new_n245_), .ZN(new_n976_));
  XOR2_X1   g775(.A(KEYINPUT127), .B(G204gat), .Z(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n974_), .B2(new_n977_), .ZN(G1353gat));
  NOR2_X1   g777(.A1(new_n971_), .A2(new_n699_), .ZN(new_n979_));
  NOR3_X1   g778(.A1(new_n979_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980_));
  XOR2_X1   g779(.A(KEYINPUT63), .B(G211gat), .Z(new_n981_));
  AOI21_X1  g780(.A(new_n980_), .B1(new_n979_), .B2(new_n981_), .ZN(G1354gat));
  OAI21_X1  g781(.A(G218gat), .B1(new_n971_), .B2(new_n687_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n697_), .A2(new_n248_), .ZN(new_n984_));
  OAI21_X1  g783(.A(new_n983_), .B1(new_n971_), .B2(new_n984_), .ZN(G1355gat));
endmodule


