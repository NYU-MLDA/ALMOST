//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT71), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT36), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G232gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT34), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n214_), .A2(new_n217_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G85gat), .B(G92gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n223_), .A2(KEYINPUT8), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(KEYINPUT8), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n228_));
  INV_X1    g027(.A(G92gat), .ZN(new_n229_));
  INV_X1    g028(.A(G85gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT64), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G85gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n229_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n228_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n217_), .A2(new_n218_), .ZN(new_n238_));
  XOR2_X1   g037(.A(KEYINPUT10), .B(G99gat), .Z(new_n239_));
  AOI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(new_n213_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n220_), .A2(new_n223_), .A3(KEYINPUT8), .A4(new_n221_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n227_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G29gat), .B(G36gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G43gat), .B(G50gat), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n249_), .A2(KEYINPUT70), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(KEYINPUT70), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n210_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n208_), .A2(new_n209_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  INV_X1    g053(.A(new_n226_), .ZN(new_n255_));
  AOI211_X1 g054(.A(new_n224_), .B(new_n255_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n256_));
  AND4_X1   g055(.A1(new_n223_), .A2(new_n220_), .A3(KEYINPUT8), .A4(new_n221_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n254_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n227_), .A2(KEYINPUT67), .A3(new_n242_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n241_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n246_), .A2(new_n247_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT15), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n246_), .A2(KEYINPUT15), .A3(new_n247_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n252_), .A2(new_n253_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n253_), .B1(new_n252_), .B2(new_n267_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n206_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n250_), .A2(new_n251_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n267_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n208_), .B(new_n209_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n252_), .A2(new_n253_), .A3(new_n267_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT36), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n205_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT72), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n270_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(KEYINPUT37), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT37), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n270_), .B(new_n278_), .C1(new_n280_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G64gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G71gat), .B(G78gat), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n286_), .A2(new_n287_), .A3(KEYINPUT11), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(KEYINPUT11), .B2(new_n286_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G1gat), .B(G8gat), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  INV_X1    g093(.A(G1gat), .ZN(new_n295_));
  INV_X1    g094(.A(G8gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n292_), .A2(new_n297_), .A3(new_n294_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n291_), .B(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G231gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G127gat), .B(G155gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G183gat), .B(G211gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT17), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n304_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n312_), .B(KEYINPUT75), .Z(new_n313_));
  AND2_X1   g112(.A1(new_n309_), .A2(new_n310_), .ZN(new_n314_));
  OR3_X1    g113(.A1(new_n304_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n285_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT76), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT22), .B(G169gat), .ZN(new_n320_));
  INV_X1    g119(.A(G176gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT82), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT80), .B(G183gat), .ZN(new_n326_));
  INV_X1    g125(.A(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G183gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT23), .B1(new_n329_), .B2(new_n327_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(G183gat), .A3(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT83), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n325_), .A2(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(KEYINPUT24), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(KEYINPUT24), .A3(new_n323_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT25), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n329_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n326_), .B2(new_n342_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT26), .B(G190gat), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n341_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n332_), .B(KEYINPUT81), .Z(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n330_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n337_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT30), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT85), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G43gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G227gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT84), .B(G15gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n352_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n351_), .A2(KEYINPUT85), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n359_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n363_), .A2(KEYINPUT86), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(KEYINPUT86), .ZN(new_n365_));
  XOR2_X1   g164(.A(G113gat), .B(G120gat), .Z(new_n366_));
  OR3_X1    g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n366_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n369_), .B(KEYINPUT31), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n362_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n359_), .B(new_n360_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n370_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G197gat), .B(G204gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT21), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G211gat), .B(G218gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G197gat), .B(G204gat), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT21), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT89), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT89), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n383_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n379_), .A2(new_n380_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT90), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n390_), .A2(KEYINPUT91), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT91), .B1(new_n390_), .B2(new_n393_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n384_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n378_), .B1(new_n396_), .B2(new_n350_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT91), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n386_), .A2(KEYINPUT89), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n381_), .A2(new_n388_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n382_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n391_), .B(KEYINPUT90), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n402_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n390_), .A2(KEYINPUT91), .A3(new_n393_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n407_), .A2(new_n408_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n348_), .B1(G183gat), .B2(G190gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n324_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n341_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT25), .B(G183gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n345_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n333_), .A3(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n409_), .A2(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n397_), .A2(new_n401_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n412_), .A2(new_n416_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n378_), .B1(new_n396_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n409_), .A2(new_n337_), .A3(new_n349_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n401_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT18), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n425_), .B(new_n426_), .Z(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n419_), .A2(new_n423_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT20), .B1(new_n409_), .B2(new_n417_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n396_), .A2(new_n350_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n400_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n397_), .A2(new_n401_), .A3(new_n418_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n427_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n377_), .B1(new_n429_), .B2(new_n434_), .ZN(new_n435_));
  OR3_X1    g234(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT2), .ZN(new_n437_));
  INV_X1    g236(.A(G141gat), .ZN(new_n438_));
  INV_X1    g237(.A(G148gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n436_), .A2(new_n440_), .A3(new_n441_), .A4(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G155gat), .A2(G162gat), .ZN(new_n444_));
  OR2_X1    g243(.A1(G155gat), .A2(G162gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(KEYINPUT1), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT1), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(G155gat), .A3(G162gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n447_), .A2(new_n449_), .A3(new_n445_), .A4(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G141gat), .B(G148gat), .Z(new_n452_));
  OAI211_X1 g251(.A(new_n451_), .B(new_n452_), .C1(new_n450_), .C2(new_n449_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n446_), .A2(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n454_), .A2(KEYINPUT29), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT28), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G228gat), .ZN(new_n458_));
  INV_X1    g257(.A(G233gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(KEYINPUT29), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n460_), .B1(new_n396_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n407_), .A2(new_n408_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n461_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT92), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT92), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n461_), .A2(new_n462_), .A3(new_n469_), .A4(new_n460_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n466_), .A2(new_n384_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n457_), .B1(new_n465_), .B2(new_n471_), .ZN(new_n472_));
  OAI22_X1  g271(.A1(new_n409_), .A2(new_n463_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n470_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n396_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n475_), .A3(new_n456_), .ZN(new_n476_));
  XOR2_X1   g275(.A(G22gat), .B(G50gat), .Z(new_n477_));
  XNOR2_X1  g276(.A(G78gat), .B(G106gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n472_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n430_), .A2(new_n431_), .A3(new_n400_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n401_), .B1(new_n397_), .B2(new_n418_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n428_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n432_), .A2(new_n433_), .A3(new_n427_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(KEYINPUT27), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n369_), .A2(new_n454_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n367_), .A2(new_n368_), .A3(new_n453_), .A4(new_n446_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT4), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT4), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n369_), .A2(new_n492_), .A3(new_n454_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n488_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G1gat), .B(G29gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(new_n230_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT0), .B(G57gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n488_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n499_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n500_));
  OR3_X1    g299(.A1(new_n494_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n498_), .B1(new_n494_), .B2(new_n500_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n435_), .A2(new_n482_), .A3(new_n487_), .A4(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n428_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT33), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n491_), .A2(new_n488_), .A3(new_n493_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n489_), .A2(new_n490_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n498_), .B1(new_n510_), .B2(new_n499_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n502_), .A2(new_n507_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n506_), .A2(new_n486_), .A3(new_n508_), .A4(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n427_), .A2(KEYINPUT32), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n432_), .A2(new_n433_), .A3(new_n514_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n503_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n482_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n505_), .B1(new_n519_), .B2(KEYINPUT94), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n521_));
  AOI211_X1 g320(.A(new_n521_), .B(new_n482_), .C1(new_n518_), .C2(new_n513_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n376_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n482_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n435_), .A2(new_n487_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n375_), .A2(new_n524_), .A3(new_n504_), .A4(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G230gat), .A2(G233gat), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n243_), .A2(new_n291_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT66), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n243_), .A2(new_n291_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n243_), .B2(new_n291_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n529_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G120gat), .B(G148gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT5), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G176gat), .B(G204gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n243_), .A2(new_n291_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n258_), .A2(new_n259_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n291_), .A2(KEYINPUT12), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n543_), .B(new_n530_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n535_), .B(new_n540_), .C1(new_n529_), .C2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT68), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n545_), .B1(new_n260_), .B2(new_n241_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n543_), .A2(new_n530_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(new_n528_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n535_), .A4(new_n540_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n548_), .A2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n552_), .A2(new_n535_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n555_), .B1(new_n556_), .B2(new_n540_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT13), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n248_), .A2(new_n301_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n262_), .A2(new_n300_), .A3(new_n299_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(G229gat), .A3(G233gat), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n264_), .A2(new_n301_), .A3(new_n265_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT77), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT79), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT78), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G169gat), .B(G197gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n570_), .B(new_n574_), .Z(new_n575_));
  NOR2_X1   g374(.A1(new_n559_), .A2(new_n575_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n319_), .A2(new_n527_), .A3(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n503_), .B(KEYINPUT96), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n295_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT38), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n279_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n270_), .A2(KEYINPUT97), .A3(new_n278_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n559_), .A2(new_n575_), .A3(new_n316_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n295_), .B1(new_n590_), .B2(new_n503_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n582_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n581_), .B2(new_n580_), .ZN(G1324gat));
  INV_X1    g392(.A(new_n525_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n577_), .A2(new_n296_), .A3(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n588_), .A2(new_n594_), .A3(new_n589_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n596_), .A2(new_n597_), .A3(G8gat), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n596_), .B2(G8gat), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n595_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT99), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(KEYINPUT99), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(G1325gat));
  INV_X1    g405(.A(G15gat), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n590_), .B2(new_n375_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT41), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n577_), .A2(new_n607_), .A3(new_n375_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1326gat));
  INV_X1    g410(.A(G22gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n482_), .B(KEYINPUT100), .Z(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n590_), .B2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n577_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1327gat));
  INV_X1    g417(.A(G29gat), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n559_), .A2(new_n575_), .A3(new_n317_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT43), .ZN(new_n621_));
  INV_X1    g420(.A(new_n285_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n527_), .B2(new_n622_), .ZN(new_n623_));
  AOI211_X1 g422(.A(KEYINPUT43), .B(new_n285_), .C1(new_n523_), .C2(new_n526_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT44), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT44), .B(new_n620_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n579_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n619_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n631_), .B1(new_n630_), .B2(new_n629_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n586_), .A2(new_n317_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n527_), .A2(new_n576_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n527_), .A2(KEYINPUT103), .A3(new_n576_), .A4(new_n633_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n619_), .A3(new_n503_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n632_), .A2(new_n639_), .ZN(G1328gat));
  NAND3_X1  g439(.A1(new_n627_), .A2(new_n594_), .A3(new_n628_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G36gat), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n525_), .A2(G36gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n636_), .A2(new_n637_), .A3(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT45), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT46), .B1(new_n646_), .B2(KEYINPUT104), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT46), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n648_), .B(new_n649_), .C1(new_n642_), .C2(new_n645_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n647_), .A2(new_n650_), .ZN(G1329gat));
  AND2_X1   g450(.A1(new_n627_), .A2(new_n628_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(G43gat), .A3(new_n375_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n638_), .A2(new_n375_), .ZN(new_n654_));
  INV_X1    g453(.A(G43gat), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n653_), .A2(KEYINPUT47), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT47), .B1(new_n653_), .B2(new_n656_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1330gat));
  AOI21_X1  g458(.A(G50gat), .B1(new_n638_), .B2(new_n613_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n482_), .A2(G50gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n652_), .B2(new_n661_), .ZN(G1331gat));
  AND4_X1   g461(.A1(new_n575_), .A2(new_n588_), .A3(new_n559_), .A4(new_n317_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(G57gat), .A3(new_n503_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT106), .ZN(new_n665_));
  INV_X1    g464(.A(G57gat), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n527_), .A2(new_n575_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n558_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n527_), .A2(KEYINPUT105), .A3(new_n575_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n319_), .A3(new_n579_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n665_), .B1(new_n666_), .B2(new_n672_), .ZN(G1332gat));
  INV_X1    g472(.A(G64gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n663_), .B2(new_n594_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT48), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n319_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n594_), .A2(new_n674_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(G1333gat));
  NAND2_X1  g478(.A1(new_n663_), .A2(new_n375_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G71gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT107), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT49), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n681_), .B(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT49), .ZN(new_n687_));
  OR3_X1    g486(.A1(new_n677_), .A2(G71gat), .A3(new_n376_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n687_), .A3(new_n688_), .ZN(G1334gat));
  INV_X1    g488(.A(G78gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n663_), .B2(new_n613_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT50), .Z(new_n692_));
  NAND2_X1  g491(.A1(new_n613_), .A2(new_n690_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n677_), .B2(new_n693_), .ZN(G1335gat));
  NAND3_X1  g493(.A1(new_n559_), .A2(new_n575_), .A3(new_n316_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT109), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n696_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n231_), .A2(new_n233_), .ZN(new_n698_));
  OR3_X1    g497(.A1(new_n697_), .A2(new_n504_), .A3(new_n698_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n669_), .A2(new_n579_), .A3(new_n633_), .A4(new_n670_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(KEYINPUT108), .A3(new_n230_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT108), .B1(new_n700_), .B2(new_n230_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1336gat));
  OAI21_X1  g505(.A(G92gat), .B1(new_n697_), .B2(new_n525_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n669_), .A2(new_n633_), .A3(new_n670_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n594_), .A2(new_n229_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(G1337gat));
  INV_X1    g509(.A(KEYINPUT111), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n375_), .A2(new_n239_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n708_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n708_), .B2(new_n712_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G99gat), .B1(new_n697_), .B2(new_n376_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1338gat));
  XNOR2_X1  g519(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n524_), .A2(G106gat), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OR3_X1    g523(.A1(new_n708_), .A2(KEYINPUT113), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT113), .B1(new_n708_), .B2(new_n724_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n696_), .B(new_n482_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G106gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G106gat), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n722_), .B1(new_n728_), .B2(new_n733_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n727_), .B(new_n721_), .C1(new_n732_), .C2(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1339gat));
  INV_X1    g535(.A(KEYINPUT13), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n557_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n557_), .A2(new_n737_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n575_), .A3(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(KEYINPUT115), .B1(new_n318_), .B2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n316_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n742_), .A2(new_n558_), .A3(new_n743_), .A4(new_n575_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n741_), .A2(KEYINPUT54), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT54), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT115), .B(new_n746_), .C1(new_n318_), .C2(new_n740_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n543_), .A2(new_n530_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n529_), .B1(new_n749_), .B2(new_n549_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT116), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(new_n546_), .B2(new_n529_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n550_), .A2(new_n551_), .A3(KEYINPUT55), .A4(new_n528_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n546_), .A2(new_n755_), .A3(new_n529_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .A4(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n539_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n575_), .B1(new_n548_), .B2(new_n554_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT56), .B1(new_n758_), .B2(KEYINPUT117), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT118), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n758_), .A2(KEYINPUT117), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT56), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n759_), .A4(new_n760_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n562_), .A2(new_n566_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n566_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n564_), .A2(new_n561_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n574_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n568_), .B2(new_n574_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n557_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n763_), .A2(new_n768_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n586_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n584_), .A2(KEYINPUT57), .A3(new_n585_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n777_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT121), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT58), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n555_), .A2(new_n775_), .A3(KEYINPUT120), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT120), .B1(new_n555_), .B2(new_n775_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n758_), .B(KEYINPUT56), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n758_), .B(new_n765_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(KEYINPUT58), .C1(new_n786_), .C2(new_n787_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n622_), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n777_), .A2(KEYINPUT121), .A3(new_n781_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n780_), .A2(new_n784_), .A3(new_n793_), .A4(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n748_), .B1(new_n795_), .B2(new_n316_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n594_), .A2(new_n482_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(new_n375_), .A3(new_n579_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(G113gat), .ZN(new_n800_));
  INV_X1    g599(.A(new_n575_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n798_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n794_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT121), .B1(new_n777_), .B2(new_n781_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n790_), .A2(new_n622_), .A3(new_n792_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n779_), .B2(new_n778_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n317_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT59), .B(new_n805_), .C1(new_n811_), .C2(new_n748_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n804_), .A2(KEYINPUT122), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT122), .B1(new_n804_), .B2(new_n812_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n575_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n802_), .B1(new_n815_), .B2(new_n800_), .ZN(G1340gat));
  INV_X1    g615(.A(G120gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n558_), .B2(KEYINPUT60), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n799_), .B(new_n818_), .C1(KEYINPUT60), .C2(new_n817_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n558_), .B1(new_n804_), .B2(new_n812_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G120gat), .B1(new_n820_), .B2(new_n821_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n819_), .B1(new_n822_), .B2(new_n823_), .ZN(G1341gat));
  INV_X1    g623(.A(G127gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n799_), .A2(new_n825_), .A3(new_n317_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n813_), .A2(new_n814_), .A3(new_n316_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n825_), .ZN(G1342gat));
  OAI211_X1 g627(.A(new_n587_), .B(new_n805_), .C1(new_n811_), .C2(new_n748_), .ZN(new_n829_));
  INV_X1    g628(.A(G134gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT124), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(KEYINPUT124), .A3(new_n830_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n813_), .A2(new_n814_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n285_), .A2(new_n830_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(G1343gat));
  INV_X1    g637(.A(new_n796_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n376_), .A2(new_n482_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n840_), .A2(new_n594_), .A3(new_n578_), .ZN(new_n841_));
  XOR2_X1   g640(.A(new_n841_), .B(KEYINPUT125), .Z(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n575_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(new_n438_), .ZN(G1344gat));
  NOR2_X1   g644(.A1(new_n843_), .A2(new_n558_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(new_n439_), .ZN(G1345gat));
  NOR2_X1   g646(.A1(new_n843_), .A2(new_n316_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT61), .B(G155gat), .Z(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  INV_X1    g649(.A(G162gat), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n843_), .A2(new_n851_), .A3(new_n285_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n843_), .B2(new_n586_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT126), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT126), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n855_), .B(new_n851_), .C1(new_n843_), .C2(new_n586_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n852_), .B1(new_n854_), .B2(new_n856_), .ZN(G1347gat));
  NAND2_X1  g656(.A1(new_n375_), .A2(new_n578_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n525_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n796_), .A2(new_n613_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G169gat), .B1(new_n862_), .B2(new_n575_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT62), .B(G169gat), .C1(new_n862_), .C2(new_n575_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n861_), .A2(new_n320_), .A3(new_n801_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(G1348gat));
  AOI21_X1  g667(.A(G176gat), .B1(new_n861_), .B2(new_n559_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n796_), .A2(new_n482_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n860_), .A2(new_n321_), .A3(new_n558_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(G1349gat));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n317_), .A3(new_n859_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n316_), .A2(new_n414_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n873_), .A2(new_n326_), .B1(new_n861_), .B2(new_n874_), .ZN(G1350gat));
  OAI21_X1  g674(.A(G190gat), .B1(new_n862_), .B2(new_n285_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n861_), .A2(new_n345_), .A3(new_n587_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1351gat));
  NOR3_X1   g677(.A1(new_n840_), .A2(new_n503_), .A3(new_n525_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n796_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n801_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n559_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g684(.A1(new_n881_), .A2(new_n317_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT63), .B(G211gat), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n886_), .B2(new_n889_), .ZN(G1354gat));
  INV_X1    g689(.A(G218gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n881_), .A2(new_n891_), .A3(new_n587_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n881_), .B2(new_n622_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT127), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n894_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(new_n892_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n895_), .A2(new_n898_), .ZN(G1355gat));
endmodule


