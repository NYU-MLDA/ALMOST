//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT85), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT1), .ZN(new_n205_));
  OR2_X1    g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n204_), .B1(new_n203_), .B2(KEYINPUT1), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT86), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n203_), .A2(KEYINPUT1), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n203_), .A2(KEYINPUT1), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT85), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT86), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(new_n206_), .A4(new_n205_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(new_n210_), .A3(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G141gat), .B(G148gat), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT87), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(KEYINPUT87), .A3(new_n216_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n206_), .A2(new_n203_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222_));
  INV_X1    g021(.A(G141gat), .ZN(new_n223_));
  INV_X1    g022(.A(G148gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(KEYINPUT88), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT88), .ZN(new_n226_));
  OAI22_X1  g025(.A1(new_n226_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(KEYINPUT89), .B2(KEYINPUT2), .ZN(new_n229_));
  AND2_X1   g028(.A1(KEYINPUT89), .A2(KEYINPUT2), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n225_), .B(new_n227_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT90), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n221_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT91), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(KEYINPUT91), .B(new_n221_), .C1(new_n231_), .C2(new_n233_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n219_), .A2(new_n220_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT28), .B1(new_n239_), .B2(KEYINPUT29), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n217_), .A2(new_n218_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT28), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .A4(new_n220_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G22gat), .B(G50gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n240_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G78gat), .B(G106gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(KEYINPUT95), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G228gat), .A2(G233gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n243_), .B1(new_n241_), .B2(new_n220_), .ZN(new_n257_));
  INV_X1    g056(.A(G197gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G204gat), .ZN(new_n259_));
  INV_X1    g058(.A(G204gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(G197gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT21), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n259_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT93), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT93), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n259_), .A2(new_n261_), .A3(new_n265_), .A4(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G211gat), .B(G218gat), .Z(new_n268_));
  INV_X1    g067(.A(KEYINPUT92), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n260_), .B2(G197gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n258_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n261_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n268_), .B1(new_n272_), .B2(KEYINPUT21), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n262_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n267_), .A2(new_n273_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n256_), .B1(new_n257_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n239_), .A2(KEYINPUT29), .ZN(new_n277_));
  INV_X1    g076(.A(new_n275_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n255_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n254_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n276_), .A2(new_n279_), .A3(new_n254_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n250_), .A2(KEYINPUT96), .A3(new_n281_), .A4(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT96), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n284_), .B1(new_n285_), .B2(new_n280_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n250_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n252_), .A2(KEYINPUT94), .ZN(new_n289_));
  INV_X1    g088(.A(new_n279_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n255_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n276_), .B(new_n279_), .C1(KEYINPUT94), .C2(new_n252_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n252_), .A2(KEYINPUT94), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n288_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n287_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT101), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT102), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n299_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G8gat), .B(G36gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT19), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT99), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT25), .B(G183gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT26), .B(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n311_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT24), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT97), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n317_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(new_n323_), .B2(new_n322_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n321_), .B(KEYINPUT98), .ZN(new_n326_));
  INV_X1    g125(.A(G169gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT22), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(G169gat), .ZN(new_n330_));
  INV_X1    g129(.A(G176gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n328_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n326_), .A2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n314_), .B(new_n315_), .C1(G183gat), .C2(G190gat), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n320_), .A2(new_n325_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n308_), .B1(new_n335_), .B2(new_n275_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n322_), .A2(new_n317_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n311_), .A2(new_n337_), .A3(new_n316_), .A4(new_n319_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n331_), .B1(new_n339_), .B2(new_n329_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G169gat), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n327_), .B(new_n331_), .C1(new_n339_), .C2(new_n329_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n334_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT20), .B1(new_n344_), .B2(new_n275_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n336_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n335_), .A2(new_n308_), .A3(new_n275_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n307_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n335_), .A2(new_n275_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n275_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n349_), .A2(KEYINPUT20), .A3(new_n350_), .A4(new_n307_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n305_), .B1(new_n348_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n335_), .A2(new_n275_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT99), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT20), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n338_), .A2(new_n343_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n278_), .B2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n358_), .A3(new_n347_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n307_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(new_n304_), .A3(new_n351_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n353_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n349_), .A2(KEYINPUT20), .A3(new_n350_), .A4(new_n360_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n345_), .B1(new_n275_), .B2(new_n335_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(new_n360_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n304_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n353_), .A2(KEYINPUT27), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n297_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G127gat), .B(G134gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G113gat), .B(G120gat), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n375_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n241_), .B2(new_n220_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n373_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n380_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n239_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n376_), .A2(new_n379_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n241_), .A2(new_n220_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(KEYINPUT4), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT105), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n385_), .A2(new_n387_), .A3(new_n373_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G1gat), .B(G29gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G85gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT0), .B(G57gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .A4(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n385_), .A2(new_n387_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n398_), .A2(new_n373_), .B1(new_n383_), .B2(new_n388_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n397_), .B1(new_n399_), .B2(new_n396_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n390_), .B1(new_n399_), .B2(new_n396_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n403_), .B(KEYINPUT82), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n357_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G71gat), .B(G99gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G15gat), .B(G43gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT81), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n344_), .A2(new_n406_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n338_), .A2(new_n343_), .A3(new_n406_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n408_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n410_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n412_), .B1(new_n410_), .B2(new_n415_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n405_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n418_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(new_n404_), .A3(new_n416_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n421_), .A3(KEYINPUT84), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n380_), .B(KEYINPUT31), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n422_), .B(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n372_), .A2(new_n402_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n371_), .B1(new_n287_), .B2(new_n296_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n385_), .A2(KEYINPUT4), .A3(new_n387_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n373_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n385_), .B2(KEYINPUT4), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n391_), .B(new_n396_), .C1(new_n428_), .C2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT103), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT33), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n385_), .A2(new_n387_), .A3(new_n429_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n395_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n381_), .A2(new_n382_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n388_), .A2(new_n373_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n437_), .B2(KEYINPUT104), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT104), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n388_), .A2(new_n439_), .A3(new_n436_), .A4(new_n373_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n363_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n431_), .A2(KEYINPUT103), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n433_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT32), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n304_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n361_), .B2(new_n351_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n446_), .B2(new_n368_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n283_), .A2(new_n286_), .B1(new_n288_), .B2(new_n295_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n402_), .A2(new_n427_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n426_), .B1(new_n452_), .B2(new_n425_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT78), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455_));
  INV_X1    g254(.A(G8gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G8gat), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n459_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G29gat), .B(G36gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G43gat), .B(G50gat), .Z(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G43gat), .B(G50gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n462_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G229gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT15), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n466_), .A2(KEYINPUT15), .A3(new_n468_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n462_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G113gat), .B(G141gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(G169gat), .B(G197gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n476_), .A2(new_n481_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n476_), .B2(new_n481_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n454_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n490_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(KEYINPUT78), .A3(new_n488_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G230gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(KEYINPUT10), .B(G99gat), .Z(new_n498_));
  INV_X1    g297(.A(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G85gat), .B(G92gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT9), .ZN(new_n502_));
  INV_X1    g301(.A(G85gat), .ZN(new_n503_));
  INV_X1    g302(.A(G92gat), .ZN(new_n504_));
  OR3_X1    g303(.A1(new_n503_), .A2(new_n504_), .A3(KEYINPUT9), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT6), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(G99gat), .A3(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n500_), .A2(new_n502_), .A3(new_n505_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512_));
  INV_X1    g311(.A(G99gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n499_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT64), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n512_), .A2(new_n513_), .A3(new_n499_), .A4(KEYINPUT64), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n516_), .A2(new_n510_), .A3(new_n517_), .A4(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT8), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT65), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n519_), .A2(new_n501_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n519_), .B2(new_n501_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n511_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G57gat), .B(G64gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT11), .ZN(new_n526_));
  XOR2_X1   g325(.A(G71gat), .B(G78gat), .Z(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n527_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n525_), .A2(KEYINPUT11), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n524_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n532_), .B(new_n511_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(KEYINPUT12), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT12), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n524_), .A2(new_n537_), .A3(new_n533_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n497_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n534_), .A2(new_n535_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n497_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G120gat), .B(G148gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT5), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G176gat), .B(G204gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n540_), .A2(new_n542_), .A3(new_n549_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n548_), .A2(KEYINPUT13), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT13), .B1(new_n548_), .B2(new_n550_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n553_), .A2(KEYINPUT66), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(KEYINPUT66), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n495_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n453_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT37), .ZN(new_n558_));
  XOR2_X1   g357(.A(G134gat), .B(G162gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT36), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT35), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n567_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n524_), .B2(new_n470_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n478_), .A2(new_n479_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n519_), .A2(new_n501_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n521_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n519_), .A2(new_n501_), .A3(new_n521_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n571_), .B1(new_n576_), .B2(new_n511_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n568_), .B1(new_n570_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n524_), .A2(new_n479_), .A3(new_n478_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n576_), .A2(new_n511_), .A3(new_n469_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n568_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .A4(new_n569_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n563_), .B1(new_n578_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n561_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT68), .B(KEYINPUT69), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n578_), .A2(new_n582_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT70), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n578_), .A2(new_n582_), .A3(KEYINPUT70), .A4(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n583_), .B1(new_n592_), .B2(KEYINPUT71), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT71), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n594_), .A3(new_n591_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n558_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n578_), .A2(new_n582_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n563_), .B1(new_n597_), .B2(KEYINPUT72), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(KEYINPUT72), .B2(new_n597_), .ZN(new_n599_));
  XOR2_X1   g398(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n592_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT74), .B1(new_n596_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n590_), .A2(new_n594_), .A3(new_n591_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n594_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n583_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n604_), .B(new_n601_), .C1(new_n607_), .C2(new_n558_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n462_), .B(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n533_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n614_), .B1(new_n617_), .B2(KEYINPUT17), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(KEYINPUT17), .B2(new_n614_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n617_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT75), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n619_), .B(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n610_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n402_), .ZN(new_n625_));
  AND4_X1   g424(.A1(new_n202_), .A2(new_n557_), .A3(new_n624_), .A4(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(KEYINPUT38), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT107), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(KEYINPUT38), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT106), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n371_), .ZN(new_n632_));
  AND4_X1   g431(.A1(new_n451_), .A2(new_n425_), .A3(new_n402_), .A4(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n450_), .A2(new_n451_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n297_), .A2(new_n402_), .A3(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n425_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n599_), .A2(new_n592_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n556_), .A2(new_n622_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n402_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n628_), .A2(new_n631_), .A3(new_n644_), .ZN(G1324gat));
  NAND3_X1  g444(.A1(new_n641_), .A2(new_n371_), .A3(new_n642_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n647_), .A3(G8gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n646_), .B2(G8gat), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n557_), .A2(new_n624_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n371_), .A2(new_n456_), .ZN(new_n652_));
  OAI22_X1  g451(.A1(new_n649_), .A2(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n643_), .B2(new_n637_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT41), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n651_), .A2(G15gat), .A3(new_n637_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1326gat));
  OAI21_X1  g458(.A(G22gat), .B1(new_n643_), .B2(new_n451_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n451_), .A2(G22gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n661_), .B1(new_n651_), .B2(new_n662_), .ZN(G1327gat));
  NOR2_X1   g462(.A1(new_n622_), .A2(new_n639_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n425_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n556_), .B(new_n664_), .C1(new_n665_), .C2(new_n633_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT110), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT110), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n453_), .A2(new_n668_), .A3(new_n556_), .A4(new_n664_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n625_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n556_), .A2(new_n623_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n603_), .A2(new_n608_), .A3(KEYINPUT108), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT43), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n610_), .C1(new_n665_), .C2(new_n633_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n676_), .B1(new_n453_), .B2(new_n610_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT44), .B(new_n674_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n676_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n638_), .B2(new_n609_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n673_), .B1(new_n682_), .B2(new_n677_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n625_), .A2(G29gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n672_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  OAI211_X1 g487(.A(new_n680_), .B(new_n371_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G36gat), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n632_), .A2(G36gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n667_), .A2(new_n669_), .A3(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n690_), .A2(KEYINPUT46), .A3(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1329gat));
  NAND2_X1  g498(.A1(new_n425_), .A2(G43gat), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n670_), .A2(new_n637_), .ZN(new_n701_));
  OAI22_X1  g500(.A1(new_n685_), .A2(new_n700_), .B1(G43gat), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g502(.A(G50gat), .B1(new_n671_), .B2(new_n297_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n297_), .A2(G50gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n686_), .B2(new_n705_), .ZN(G1331gat));
  NAND2_X1  g505(.A1(new_n554_), .A2(new_n555_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n622_), .A2(new_n495_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n641_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(G57gat), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n402_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT114), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n610_), .A2(new_n707_), .A3(new_n623_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n714_), .A2(KEYINPUT112), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n638_), .A2(new_n494_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n707_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n624_), .A2(KEYINPUT112), .A3(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n715_), .A2(new_n716_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n715_), .A2(new_n716_), .A3(KEYINPUT113), .A4(new_n718_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n625_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n713_), .B1(new_n711_), .B2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(KEYINPUT115), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n632_), .A2(G64gat), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n721_), .A2(new_n722_), .A3(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G64gat), .B1(new_n710_), .B2(new_n632_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n725_), .B1(new_n727_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n728_), .B(KEYINPUT48), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n721_), .A2(new_n722_), .A3(new_n726_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(KEYINPUT115), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n710_), .B2(new_n637_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT49), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n637_), .A2(G71gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n721_), .A2(new_n722_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n710_), .B2(new_n451_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n451_), .A2(G78gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n721_), .A2(new_n722_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1335gat));
  NAND2_X1  g544(.A1(new_n682_), .A2(new_n677_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n717_), .A2(new_n623_), .A3(new_n495_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n402_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n707_), .A2(new_n639_), .A3(new_n622_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n716_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n503_), .A3(new_n625_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n750_), .A2(new_n754_), .ZN(G1336gat));
  OAI21_X1  g554(.A(G92gat), .B1(new_n749_), .B2(new_n632_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(new_n504_), .A3(new_n371_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n749_), .B2(new_n637_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n753_), .A2(new_n498_), .A3(new_n425_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g561(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n763_));
  AOI211_X1 g562(.A(new_n451_), .B(new_n747_), .C1(new_n682_), .C2(new_n677_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT52), .B1(new_n764_), .B2(new_n499_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n746_), .A2(new_n297_), .A3(new_n748_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n765_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n297_), .A2(new_n499_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n752_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n763_), .B1(new_n769_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n763_), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n771_), .B(new_n774_), .C1(new_n765_), .C2(new_n768_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n536_), .A2(new_n497_), .A3(new_n538_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n778_), .A2(new_n539_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n536_), .A2(new_n538_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n779_), .A3(new_n496_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n547_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n777_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n549_), .B1(new_n539_), .B2(new_n779_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n540_), .A2(KEYINPUT55), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT56), .B(new_n785_), .C1(new_n786_), .C2(new_n778_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n550_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n473_), .A2(new_n474_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n480_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n486_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n488_), .A2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT117), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n789_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n788_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n788_), .A2(KEYINPUT58), .A3(new_n795_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n603_), .A2(new_n608_), .A3(new_n798_), .A4(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n494_), .A2(new_n550_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n794_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n639_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n800_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT57), .B1(new_n804_), .B2(KEYINPUT118), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n809_), .B(new_n639_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n807_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n623_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n708_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n609_), .A2(new_n814_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n815_), .A2(KEYINPUT54), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(KEYINPUT54), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n813_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n372_), .A2(new_n625_), .A3(new_n425_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n820_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n804_), .A2(KEYINPUT118), .ZN(new_n825_));
  AND4_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n805_), .A4(new_n810_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n824_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n807_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT120), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n807_), .B(new_n830_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n623_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n821_), .B1(new_n832_), .B2(new_n818_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n494_), .B(new_n823_), .C1(new_n833_), .C2(new_n820_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G113gat), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n818_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n822_), .ZN(new_n837_));
  OR3_X1    g636(.A1(new_n837_), .A2(G113gat), .A3(new_n495_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(G1340gat));
  OAI211_X1 g638(.A(new_n717_), .B(new_n823_), .C1(new_n833_), .C2(new_n820_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G120gat), .ZN(new_n841_));
  INV_X1    g640(.A(G120gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n707_), .B2(KEYINPUT60), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n833_), .B(new_n843_), .C1(KEYINPUT60), .C2(new_n842_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(G1341gat));
  AOI21_X1  g644(.A(G127gat), .B1(new_n833_), .B2(new_n622_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n823_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n837_), .B2(KEYINPUT59), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n622_), .A2(G127gat), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(KEYINPUT121), .Z(new_n850_));
  AOI21_X1  g649(.A(new_n846_), .B1(new_n848_), .B2(new_n850_), .ZN(G1342gat));
  OAI211_X1 g650(.A(new_n610_), .B(new_n823_), .C1(new_n833_), .C2(new_n820_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G134gat), .ZN(new_n853_));
  OR3_X1    g652(.A1(new_n837_), .A2(G134gat), .A3(new_n639_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1343gat));
  AOI21_X1  g654(.A(new_n425_), .B1(new_n832_), .B2(new_n818_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n451_), .A2(new_n402_), .A3(new_n371_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n494_), .A3(new_n857_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT122), .B(G141gat), .Z(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1344gat));
  NAND3_X1  g659(.A1(new_n856_), .A2(new_n717_), .A3(new_n857_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT123), .B(G148gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1345gat));
  NAND3_X1  g662(.A1(new_n856_), .A2(new_n622_), .A3(new_n857_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  INV_X1    g665(.A(G162gat), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n856_), .A2(new_n867_), .A3(new_n640_), .A4(new_n857_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n856_), .A2(new_n610_), .A3(new_n857_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n625_), .A2(new_n632_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n425_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n819_), .A2(new_n451_), .A3(new_n494_), .A4(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT124), .B1(new_n874_), .B2(G169gat), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(KEYINPUT62), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n328_), .A2(new_n330_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n874_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n875_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n882_), .ZN(G1348gat));
  NAND2_X1  g682(.A1(new_n819_), .A2(new_n451_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n872_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G176gat), .B1(new_n885_), .B2(new_n717_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n297_), .B1(new_n832_), .B2(new_n818_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n707_), .A2(new_n331_), .A3(new_n872_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1349gat));
  NOR2_X1   g688(.A1(new_n872_), .A2(new_n623_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G183gat), .B1(new_n887_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n890_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n884_), .A2(new_n309_), .A3(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT125), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  OR3_X1    g693(.A1(new_n884_), .A2(new_n309_), .A3(new_n892_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896_));
  AOI211_X1 g695(.A(new_n297_), .B(new_n892_), .C1(new_n832_), .C2(new_n818_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n895_), .B(new_n896_), .C1(new_n897_), .C2(G183gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n898_), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n885_), .A2(new_n640_), .A3(new_n310_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n884_), .A2(new_n609_), .A3(new_n872_), .ZN(new_n901_));
  INV_X1    g700(.A(G190gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1351gat));
  NOR3_X1   g702(.A1(new_n451_), .A2(new_n625_), .A3(new_n632_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n856_), .A2(new_n494_), .A3(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT126), .B(G197gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1352gat));
  NAND3_X1  g706(.A1(new_n856_), .A2(new_n717_), .A3(new_n904_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g708(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n836_), .A2(new_n637_), .A3(new_n904_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n623_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n913_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n856_), .A2(new_n904_), .A3(new_n915_), .A4(new_n911_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1354gat));
  OAI21_X1  g718(.A(G218gat), .B1(new_n914_), .B2(new_n609_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n639_), .A2(G218gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n914_), .B2(new_n921_), .ZN(G1355gat));
endmodule


