//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G15gat), .B(G22gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT72), .B(G8gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G1gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n208_), .B2(KEYINPUT14), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT73), .Z(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n209_), .B(KEYINPUT73), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(new_n211_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G29gat), .B(G36gat), .Z(new_n217_));
  XOR2_X1   g016(.A(G43gat), .B(G50gat), .Z(new_n218_));
  XOR2_X1   g017(.A(new_n217_), .B(new_n218_), .Z(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n222_), .B(KEYINPUT78), .Z(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n219_), .B(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n213_), .A2(new_n226_), .A3(new_n215_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT77), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n213_), .A2(new_n215_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT77), .A3(new_n226_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n224_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n219_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n222_), .B1(new_n233_), .B2(new_n221_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n205_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n221_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n222_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n231_), .A2(new_n229_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n238_), .B(new_n204_), .C1(new_n239_), .C2(new_n224_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT23), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(G183gat), .A3(G190gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT24), .ZN(new_n247_));
  NOR2_X1   g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n244_), .A2(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(KEYINPUT24), .A3(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT25), .B(G183gat), .ZN(new_n257_));
  INV_X1    g056(.A(G190gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT26), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT79), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G190gat), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n257_), .B(new_n261_), .C1(new_n262_), .C2(new_n260_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT80), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT26), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(G190gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n259_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT79), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n269_), .A2(KEYINPUT80), .A3(new_n257_), .A4(new_n261_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n256_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT22), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G169gat), .ZN(new_n274_));
  INV_X1    g073(.A(G169gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT22), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT82), .ZN(new_n278_));
  OR2_X1    g077(.A1(KEYINPUT83), .A2(G176gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(KEYINPUT83), .A2(G176gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT82), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n274_), .A2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n278_), .A2(new_n282_), .A3(KEYINPUT84), .A4(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT84), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n275_), .A2(KEYINPUT22), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n279_), .B(new_n280_), .C1(new_n287_), .C2(KEYINPUT82), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n286_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n244_), .A2(new_n246_), .A3(KEYINPUT85), .ZN(new_n292_));
  INV_X1    g091(.A(G183gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n258_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n295_), .A2(new_n245_), .A3(G183gat), .A4(G190gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n297_), .A2(new_n253_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n291_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n272_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G71gat), .B(G99gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n301_), .B(G43gat), .Z(new_n302_));
  NOR2_X1   g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n256_), .A2(new_n271_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n302_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n307_));
  OR3_X1    g106(.A1(new_n303_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n307_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G127gat), .B(G134gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G113gat), .B(G120gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n313_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(KEYINPUT86), .A3(new_n316_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(G15gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT30), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n321_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n310_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT88), .ZN(new_n328_));
  AND2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT92), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335_));
  INV_X1    g134(.A(G141gat), .ZN(new_n336_));
  INV_X1    g135(.A(G148gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n332_), .B1(new_n334_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT91), .ZN(new_n344_));
  OR2_X1    g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n345_), .B1(KEYINPUT1), .B2(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n346_), .A2(KEYINPUT90), .A3(KEYINPUT1), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT90), .B1(new_n346_), .B2(KEYINPUT1), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT89), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(G141gat), .B2(G148gat), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n351_), .A2(new_n353_), .B1(G141gat), .B2(G148gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n344_), .B1(new_n350_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT1), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n330_), .B1(new_n329_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n346_), .A2(KEYINPUT1), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT90), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n346_), .A2(KEYINPUT90), .A3(KEYINPUT1), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT91), .A3(new_n354_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n343_), .B1(new_n356_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n367_), .A2(KEYINPUT28), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(KEYINPUT28), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G197gat), .A2(G204gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G197gat), .A2(G204gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT94), .ZN(new_n375_));
  INV_X1    g174(.A(G211gat), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(KEYINPUT21), .A4(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n378_), .A2(new_n375_), .A3(KEYINPUT21), .A4(new_n371_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G211gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G218gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n371_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT21), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n372_), .A2(new_n373_), .A3(new_n384_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT93), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(KEYINPUT93), .A3(new_n384_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n381_), .A2(new_n382_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n377_), .A2(new_n380_), .A3(G218gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n333_), .B(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n331_), .B1(new_n394_), .B2(new_n341_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n363_), .A2(KEYINPUT91), .A3(new_n354_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT91), .B1(new_n363_), .B2(new_n354_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n392_), .B1(new_n398_), .B2(KEYINPUT29), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n370_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(G78gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G106gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G22gat), .B(G50gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n403_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n400_), .A2(new_n402_), .A3(new_n410_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT18), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT32), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n304_), .B2(new_n392_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n381_), .A2(new_n382_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n388_), .A2(new_n389_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n424_), .A2(new_n391_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n248_), .A2(new_n247_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n257_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n254_), .B(new_n427_), .C1(new_n428_), .C2(new_n268_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n292_), .A2(new_n296_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n253_), .B1(new_n281_), .B2(new_n277_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n244_), .A2(new_n246_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n432_), .A2(new_n294_), .ZN(new_n433_));
  OAI22_X1  g232(.A1(new_n429_), .A2(new_n430_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n426_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n423_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G226gat), .A2(G233gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT19), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n422_), .B1(new_n300_), .B2(new_n426_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n434_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n440_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n421_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n436_), .A2(new_n438_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n441_), .A2(new_n443_), .A3(new_n440_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(new_n420_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G1gat), .B(G29gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n317_), .B(new_n395_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n315_), .A2(KEYINPUT86), .A3(new_n316_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT86), .B1(new_n315_), .B2(new_n316_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n455_), .B1(new_n365_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G225gat), .A2(G233gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n454_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n455_), .B(KEYINPUT4), .C1(new_n365_), .C2(new_n458_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n463_), .A2(new_n461_), .ZN(new_n464_));
  XOR2_X1   g263(.A(KEYINPUT95), .B(KEYINPUT4), .Z(new_n465_));
  NAND3_X1  g264(.A1(new_n398_), .A2(new_n321_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT96), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n398_), .A2(new_n321_), .A3(KEYINPUT96), .A4(new_n465_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n462_), .B1(new_n464_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n454_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n463_), .A2(new_n461_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n474_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n459_), .A2(new_n461_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n473_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n449_), .B1(new_n472_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT98), .B1(new_n471_), .B2(KEYINPUT33), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT98), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n481_), .B(new_n482_), .C1(new_n475_), .C2(new_n462_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT99), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n459_), .A2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n455_), .B(KEYINPUT99), .C1(new_n365_), .C2(new_n458_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n461_), .A3(new_n487_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n468_), .A2(new_n469_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n463_), .A2(new_n460_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n488_), .B(new_n473_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT20), .B1(new_n304_), .B2(new_n392_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n492_), .A2(new_n438_), .A3(new_n442_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n440_), .B1(new_n423_), .B2(new_n435_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n418_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n446_), .A2(new_n447_), .A3(new_n419_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n491_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n471_), .A2(KEYINPUT33), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n484_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n479_), .B1(new_n499_), .B2(KEYINPUT100), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT100), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n484_), .A2(new_n497_), .A3(new_n501_), .A4(new_n498_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n414_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n478_), .A2(new_n472_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n496_), .A2(new_n495_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT27), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n418_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(KEYINPUT27), .A3(new_n496_), .ZN(new_n510_));
  AND4_X1   g309(.A1(new_n505_), .A2(new_n414_), .A3(new_n508_), .A4(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n328_), .B1(new_n503_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n414_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n327_), .A2(new_n505_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT101), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT101), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n508_), .A2(new_n510_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n513_), .A4(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n242_), .B1(new_n512_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT37), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT65), .ZN(new_n525_));
  OR3_X1    g324(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n528_), .A2(KEYINPUT66), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT6), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n525_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  OR3_X1    g332(.A1(new_n532_), .A2(KEYINPUT66), .A3(new_n528_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G85gat), .B(G92gat), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n524_), .B1(new_n538_), .B2(KEYINPUT65), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(G85gat), .ZN(new_n541_));
  INV_X1    g340(.A(G92gat), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n541_), .A2(new_n542_), .A3(KEYINPUT9), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT10), .B(G99gat), .Z(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n544_), .B2(new_n407_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n536_), .A2(KEYINPUT9), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(KEYINPUT8), .B2(new_n528_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n540_), .B1(new_n548_), .B2(new_n531_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n537_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(new_n219_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n551_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n226_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(KEYINPUT71), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n555_), .A2(new_n552_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n565_));
  INV_X1    g364(.A(new_n560_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n556_), .B(new_n557_), .C1(KEYINPUT71), .C2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n561_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n561_), .A2(new_n567_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n564_), .B(KEYINPUT36), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n523_), .B(new_n568_), .C1(new_n569_), .C2(new_n571_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n561_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n571_), .B1(new_n561_), .B2(new_n567_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT37), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT11), .ZN(new_n578_));
  XOR2_X1   g377(.A(G71gat), .B(G78gat), .Z(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n577_), .A2(KEYINPUT11), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n580_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n216_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT75), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n216_), .A2(new_n586_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G127gat), .B(G155gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n590_), .B(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n587_), .A2(new_n589_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(new_n596_), .A3(new_n595_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT76), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n576_), .A2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G120gat), .B(G148gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(G176gat), .B(G204gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT68), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT64), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n584_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n537_), .A2(new_n549_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n538_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n528_), .A2(KEYINPUT8), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n546_), .B2(new_n545_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n539_), .B1(new_n617_), .B2(new_n532_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n584_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(new_n619_), .A3(KEYINPUT12), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT12), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n550_), .A2(new_n621_), .A3(new_n584_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n612_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n611_), .B1(new_n614_), .B2(new_n619_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n609_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n623_), .A2(new_n624_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT69), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n608_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n626_), .B2(new_n608_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n625_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT13), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n608_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT69), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n628_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(KEYINPUT13), .A3(new_n625_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n603_), .A2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n522_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(G1gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n504_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT38), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n573_), .A2(new_n574_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n512_), .B2(new_n521_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n601_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n638_), .A2(new_n646_), .A3(new_n242_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(KEYINPUT102), .A3(new_n647_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n505_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n641_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n652_), .A2(KEYINPUT103), .A3(new_n641_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n643_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(KEYINPUT104), .B(new_n643_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1324gat));
  INV_X1    g460(.A(new_n519_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n645_), .A2(new_n662_), .A3(new_n647_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT105), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G8gat), .B1(new_n663_), .B2(KEYINPUT105), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT106), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT39), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n663_), .A2(KEYINPUT105), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(G8gat), .A4(new_n664_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n667_), .A2(new_n671_), .A3(KEYINPUT39), .ZN(new_n672_));
  INV_X1    g471(.A(new_n207_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n640_), .A2(new_n662_), .A3(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n668_), .A2(new_n672_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n668_), .A2(KEYINPUT40), .A3(new_n672_), .A4(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  INV_X1    g478(.A(G15gat), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n650_), .A2(new_n651_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n328_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n680_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT41), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n640_), .A2(new_n680_), .A3(new_n682_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1326gat));
  INV_X1    g485(.A(G22gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n681_), .B2(new_n414_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT42), .Z(new_n689_));
  NAND3_X1  g488(.A1(new_n640_), .A2(new_n687_), .A3(new_n414_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1327gat));
  NOR3_X1   g490(.A1(new_n602_), .A2(new_n638_), .A3(new_n242_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n480_), .A2(new_n483_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n498_), .A2(new_n496_), .A3(new_n495_), .A4(new_n491_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT100), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n504_), .A2(new_n445_), .A3(new_n448_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n502_), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n511_), .B1(new_n697_), .B2(new_n513_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n521_), .B1(new_n698_), .B2(new_n682_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n576_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n699_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n692_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n697_), .A2(new_n513_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n511_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n682_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n516_), .A2(new_n520_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n700_), .B(new_n701_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n576_), .B1(new_n512_), .B2(new_n521_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n703_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(KEYINPUT44), .A3(new_n692_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n707_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n504_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G29gat), .ZN(new_n718_));
  INV_X1    g517(.A(new_n644_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n602_), .A2(new_n638_), .A3(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n522_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n505_), .A2(G29gat), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT108), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n718_), .B1(new_n722_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g524(.A(G36gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n716_), .B2(new_n662_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n721_), .A2(new_n726_), .A3(new_n662_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT45), .Z(new_n729_));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  OR3_X1    g529(.A1(new_n727_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1329gat));
  AND2_X1   g532(.A1(new_n327_), .A2(G43gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n716_), .A2(KEYINPUT109), .A3(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT110), .B(G43gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n722_), .B2(new_n328_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n707_), .A2(new_n715_), .A3(new_n734_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n737_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT47), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n735_), .A2(new_n743_), .A3(new_n737_), .A4(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1330gat));
  AOI21_X1  g544(.A(G50gat), .B1(new_n721_), .B2(new_n414_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n414_), .A2(G50gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n716_), .B2(new_n747_), .ZN(G1331gat));
  INV_X1    g547(.A(new_n638_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n241_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n645_), .A2(new_n602_), .A3(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(G57gat), .A3(new_n504_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(KEYINPUT111), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(KEYINPUT111), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n699_), .A2(new_n750_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n602_), .A3(new_n576_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G57gat), .B1(new_n757_), .B2(new_n504_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n753_), .A2(new_n754_), .A3(new_n758_), .ZN(G1332gat));
  INV_X1    g558(.A(G64gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n751_), .B2(new_n662_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n757_), .A2(new_n760_), .A3(new_n662_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1333gat));
  INV_X1    g564(.A(G71gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n751_), .B2(new_n682_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT49), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n757_), .A2(new_n766_), .A3(new_n682_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1334gat));
  AOI21_X1  g569(.A(new_n405_), .B1(new_n751_), .B2(new_n414_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT50), .Z(new_n772_));
  NAND2_X1  g571(.A1(new_n414_), .A2(new_n405_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT113), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n772_), .B1(new_n756_), .B2(new_n774_), .ZN(G1335gat));
  INV_X1    g574(.A(new_n755_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n776_), .A2(new_n719_), .A3(new_n602_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(new_n541_), .A3(new_n504_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n750_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n779_), .A2(new_n602_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n714_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n504_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n778_), .B1(new_n783_), .B2(new_n541_), .ZN(G1336gat));
  NAND3_X1  g583(.A1(new_n777_), .A2(new_n542_), .A3(new_n662_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n781_), .A2(new_n662_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n787_), .B2(new_n542_), .ZN(G1337gat));
  OAI211_X1 g587(.A(new_n682_), .B(new_n780_), .C1(new_n702_), .C2(new_n704_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(G99gat), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT114), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n792_), .A2(KEYINPUT51), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n327_), .A2(new_n544_), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n777_), .A2(new_n794_), .B1(new_n792_), .B2(KEYINPUT51), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n793_), .B1(new_n791_), .B2(new_n795_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n777_), .A2(new_n407_), .A3(new_n414_), .ZN(new_n800_));
  XOR2_X1   g599(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n714_), .A2(new_n802_), .A3(new_n414_), .A4(new_n780_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(G106gat), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n414_), .B(new_n780_), .C1(new_n702_), .C2(new_n704_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT116), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n801_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  AND4_X1   g606(.A1(G106gat), .A2(new_n806_), .A3(new_n803_), .A4(new_n801_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n800_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT53), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n800_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1339gat));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n639_), .A2(new_n814_), .A3(new_n242_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n749_), .A2(new_n242_), .A3(new_n602_), .A4(new_n576_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT54), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n236_), .A2(new_n223_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n223_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n221_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n820_), .B(new_n205_), .C1(new_n239_), .C2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n823_), .A2(new_n240_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n620_), .A2(new_n612_), .A3(new_n622_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n623_), .A2(KEYINPUT55), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n623_), .B1(KEYINPUT55), .B2(new_n825_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n609_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n824_), .B(new_n636_), .C1(KEYINPUT56), .C2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(KEYINPUT56), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n819_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n824_), .A2(new_n636_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n828_), .A2(KEYINPUT56), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n830_), .A4(new_n834_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n832_), .A2(new_n700_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n828_), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n838_));
  NOR2_X1   g637(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n609_), .B(new_n839_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n838_), .A2(new_n241_), .A3(new_n636_), .A4(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n631_), .A2(new_n824_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n644_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n837_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n636_), .A2(new_n241_), .A3(new_n840_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n846_), .A2(new_n838_), .B1(new_n631_), .B2(new_n824_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT119), .B(KEYINPUT57), .C1(new_n847_), .C2(new_n644_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n836_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n818_), .B1(new_n849_), .B2(new_n602_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n327_), .A2(new_n504_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n514_), .A2(KEYINPUT59), .A3(new_n852_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n850_), .A2(new_n851_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n851_), .B1(new_n850_), .B2(new_n853_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n848_), .A2(new_n845_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n836_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n601_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n816_), .B(new_n814_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT120), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n514_), .A2(new_n852_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n818_), .B(new_n863_), .C1(new_n849_), .C2(new_n601_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n862_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT59), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n856_), .A2(new_n866_), .A3(new_n241_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(G113gat), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n242_), .A2(G113gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n865_), .B2(new_n869_), .ZN(G1340gat));
  NAND3_X1  g669(.A1(new_n856_), .A2(new_n866_), .A3(new_n638_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G120gat), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n873_));
  AOI21_X1  g672(.A(G120gat), .B1(new_n638_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT122), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n873_), .B2(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n872_), .B1(new_n865_), .B2(new_n878_), .ZN(G1341gat));
  AND3_X1   g678(.A1(new_n856_), .A2(new_n866_), .A3(new_n601_), .ZN(new_n880_));
  INV_X1    g679(.A(G127gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n602_), .A2(new_n881_), .ZN(new_n882_));
  OAI22_X1  g681(.A1(new_n880_), .A2(new_n881_), .B1(new_n865_), .B2(new_n882_), .ZN(G1342gat));
  NAND3_X1  g682(.A1(new_n856_), .A2(new_n866_), .A3(new_n700_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G134gat), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n719_), .A2(G134gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n865_), .B2(new_n886_), .ZN(G1343gat));
  AND2_X1   g686(.A1(new_n861_), .A2(new_n864_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n682_), .A2(new_n662_), .A3(new_n505_), .A4(new_n513_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n241_), .A3(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g690(.A1(new_n888_), .A2(new_n638_), .A3(new_n889_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g692(.A1(new_n888_), .A2(new_n602_), .A3(new_n889_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  NAND4_X1  g695(.A1(new_n861_), .A2(new_n644_), .A3(new_n864_), .A4(new_n889_), .ZN(new_n897_));
  INV_X1    g696(.A(G162gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n899_), .A2(KEYINPUT123), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(KEYINPUT123), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n888_), .A2(new_n889_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n576_), .A2(new_n898_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n900_), .A2(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1347gat));
  INV_X1    g703(.A(new_n850_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n662_), .A2(new_n505_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n328_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n414_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n905_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n242_), .A2(new_n277_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT124), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n911_), .A2(new_n241_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(G169gat), .ZN(new_n917_));
  AOI211_X1 g716(.A(KEYINPUT62), .B(new_n275_), .C1(new_n911_), .C2(new_n241_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n914_), .B1(new_n917_), .B2(new_n918_), .ZN(G1348gat));
  AOI21_X1  g718(.A(new_n281_), .B1(new_n911_), .B2(new_n638_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n861_), .A2(new_n864_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n414_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n861_), .A2(KEYINPUT125), .A3(new_n513_), .A4(new_n864_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n907_), .A2(G176gat), .A3(new_n638_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n920_), .B1(new_n925_), .B2(new_n926_), .ZN(G1349gat));
  NAND4_X1  g726(.A1(new_n850_), .A2(new_n428_), .A3(new_n601_), .A4(new_n909_), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT126), .Z(new_n929_));
  AND2_X1   g728(.A1(new_n907_), .A2(new_n602_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n925_), .A2(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n931_), .B2(new_n293_), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n911_), .A2(new_n644_), .A3(new_n262_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n905_), .A2(new_n576_), .A3(new_n910_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n258_), .B2(new_n934_), .ZN(G1351gat));
  NOR3_X1   g734(.A1(new_n682_), .A2(new_n906_), .A3(new_n513_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n888_), .A2(new_n241_), .A3(new_n936_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g737(.A1(new_n888_), .A2(new_n638_), .A3(new_n936_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g739(.A(new_n646_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n861_), .A2(new_n864_), .A3(new_n936_), .A4(new_n941_), .ZN(new_n942_));
  AND2_X1   g741(.A1(new_n942_), .A2(KEYINPUT127), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n942_), .A2(KEYINPUT127), .ZN(new_n944_));
  NOR2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n943_), .A2(new_n944_), .A3(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n888_), .A2(new_n948_), .A3(new_n936_), .A4(new_n941_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n942_), .A2(KEYINPUT127), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n945_), .B1(new_n949_), .B2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n947_), .A2(new_n951_), .ZN(G1354gat));
  NAND2_X1  g751(.A1(new_n888_), .A2(new_n936_), .ZN(new_n953_));
  OAI21_X1  g752(.A(G218gat), .B1(new_n953_), .B2(new_n576_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n644_), .A2(new_n382_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n953_), .B2(new_n955_), .ZN(G1355gat));
endmodule


