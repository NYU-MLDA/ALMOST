//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT4), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT89), .B(G113gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G120gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(G127gat), .B(G134gat), .Z(new_n207_));
  OR2_X1    g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n207_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n219_), .B1(new_n213_), .B2(KEYINPUT1), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT92), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(KEYINPUT92), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n219_), .B(KEYINPUT3), .ZN(new_n225_));
  NAND2_X1  g024(.A1(KEYINPUT93), .A2(KEYINPUT2), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT93), .A2(KEYINPUT2), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(new_n218_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n225_), .B(new_n228_), .C1(new_n218_), .C2(new_n226_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n215_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n208_), .A2(KEYINPUT90), .A3(new_n209_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n212_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n222_), .A2(new_n223_), .B1(new_n215_), .B2(new_n229_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n210_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n204_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n208_), .A2(KEYINPUT90), .A3(new_n209_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT90), .B1(new_n208_), .B2(new_n209_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT4), .B1(new_n239_), .B2(new_n231_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n203_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT103), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n233_), .A2(new_n242_), .A3(new_n202_), .A4(new_n235_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n233_), .A2(new_n235_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT103), .B1(new_n244_), .B2(new_n203_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT0), .B(G57gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(G85gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(G1gat), .B(G29gat), .Z(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT106), .ZN(new_n252_));
  INV_X1    g051(.A(new_n250_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n241_), .A2(new_n243_), .A3(new_n245_), .A4(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n246_), .A2(KEYINPUT106), .A3(new_n250_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT18), .B(G64gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(G92gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G8gat), .B(G36gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT102), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT98), .ZN(new_n265_));
  INV_X1    g064(.A(G197gat), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n266_), .A2(G204gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(G204gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n265_), .B1(KEYINPUT21), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT97), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT96), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n268_), .B(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n267_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n271_), .B1(new_n274_), .B2(KEYINPUT21), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT21), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n273_), .A2(KEYINPUT97), .A3(new_n276_), .A4(new_n267_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n270_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n265_), .A2(new_n274_), .A3(KEYINPUT21), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT23), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT88), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n288_), .B2(KEYINPUT24), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT26), .B(G190gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT87), .ZN(new_n293_));
  INV_X1    g092(.A(G183gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n293_), .B1(new_n294_), .B2(KEYINPUT25), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT25), .B(G183gat), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n292_), .B(new_n295_), .C1(new_n296_), .C2(new_n293_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n289_), .A2(new_n291_), .A3(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n282_), .B1(G183gat), .B2(G190gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT22), .B(G169gat), .ZN(new_n300_));
  INV_X1    g099(.A(G176gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n287_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n263_), .B1(new_n280_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT101), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n286_), .A2(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n299_), .B(new_n308_), .C1(new_n307_), .C2(new_n302_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n284_), .A2(new_n290_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n296_), .A2(new_n292_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n289_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n280_), .A2(new_n309_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n278_), .A2(new_n279_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(KEYINPUT102), .A3(new_n304_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n306_), .A2(new_n313_), .A3(KEYINPUT20), .A4(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT100), .Z(new_n318_));
  XOR2_X1   g117(.A(new_n318_), .B(KEYINPUT19), .Z(new_n319_));
  AND2_X1   g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT20), .B1(new_n314_), .B2(new_n304_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n278_), .A2(new_n279_), .B1(new_n312_), .B2(new_n309_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n321_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n262_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n319_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n316_), .A2(new_n325_), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n321_), .A2(new_n325_), .A3(new_n322_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n261_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n330_), .A3(KEYINPUT27), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT27), .ZN(new_n332_));
  AOI211_X1 g131(.A(new_n261_), .B(new_n327_), .C1(new_n316_), .C2(new_n325_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n262_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT95), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n314_), .B(new_n337_), .C1(new_n338_), .C2(new_n234_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT99), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G228gat), .A2(G233gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n342_), .B(KEYINPUT94), .Z(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n314_), .B(KEYINPUT99), .C1(new_n338_), .C2(new_n234_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n339_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G22gat), .B(G50gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(G78gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n346_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n352_));
  INV_X1    g151(.A(G106gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n234_), .A2(new_n338_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n354_), .A2(KEYINPUT28), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(KEYINPUT28), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n353_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n355_), .A2(new_n353_), .A3(new_n356_), .ZN(new_n358_));
  OAI22_X1  g157(.A1(new_n351_), .A2(new_n352_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n346_), .A2(new_n347_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n349_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n358_), .A2(new_n357_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n346_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT30), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n239_), .A2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT30), .B1(new_n237_), .B2(new_n238_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n304_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n369_), .A3(new_n305_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G15gat), .B(G43gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT31), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G71gat), .B(G99gat), .Z(new_n377_));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n375_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n371_), .A2(new_n372_), .A3(new_n380_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n376_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n379_), .B1(new_n376_), .B2(new_n381_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AND4_X1   g183(.A1(new_n257_), .A2(new_n336_), .A3(new_n366_), .A4(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n333_), .A2(new_n334_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n254_), .A2(KEYINPUT104), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT33), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n202_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n244_), .B(KEYINPUT105), .Z(new_n390_));
  OAI211_X1 g189(.A(new_n250_), .B(new_n389_), .C1(new_n390_), .C2(new_n202_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT33), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n254_), .A2(KEYINPUT104), .A3(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n386_), .A2(new_n388_), .A3(new_n391_), .A4(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(KEYINPUT32), .B(new_n261_), .C1(new_n320_), .C2(new_n323_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT32), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n329_), .B1(new_n396_), .B2(new_n262_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n255_), .A2(new_n256_), .A3(new_n395_), .A4(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n394_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n366_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n336_), .A2(KEYINPUT107), .A3(new_n257_), .A4(new_n365_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n257_), .A2(new_n365_), .A3(new_n335_), .A4(new_n331_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT107), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n384_), .B(KEYINPUT91), .Z(new_n406_));
  AOI21_X1  g205(.A(new_n385_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(G1gat), .ZN(new_n408_));
  INV_X1    g207(.A(G8gat), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT14), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT78), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT78), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n412_), .B(KEYINPUT14), .C1(new_n408_), .C2(new_n409_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G15gat), .B(G22gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT79), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G1gat), .B(G8gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G231gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT80), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n418_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G71gat), .ZN(new_n422_));
  INV_X1    g221(.A(G78gat), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n423_), .A2(KEYINPUT70), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(KEYINPUT70), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n422_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT70), .B(G78gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(G71gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G57gat), .A2(G64gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT11), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G57gat), .A2(G64gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n426_), .A2(new_n428_), .A3(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(G57gat), .A2(G64gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT11), .B1(new_n435_), .B2(new_n429_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT71), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT71), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n438_), .B(KEYINPUT11), .C1(new_n435_), .C2(new_n429_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n434_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n434_), .A2(new_n440_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n421_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(G155gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G183gat), .B(G211gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT82), .B(G127gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n448_), .B(new_n449_), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT17), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n444_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n444_), .A2(KEYINPUT17), .A3(new_n450_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n407_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G230gat), .ZN(new_n456_));
  INV_X1    g255(.A(G233gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n441_), .A2(new_n442_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G99gat), .A2(G106gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT67), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n461_), .A2(KEYINPUT6), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(KEYINPUT67), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(KEYINPUT67), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(KEYINPUT6), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n466_), .A2(new_n467_), .A3(G99gat), .A4(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n469_));
  INV_X1    g268(.A(G99gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n353_), .ZN(new_n471_));
  AND2_X1   g270(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n472_));
  NOR2_X1   g271(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n473_));
  OAI22_X1  g272(.A1(new_n472_), .A2(new_n473_), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n465_), .A2(new_n468_), .A3(new_n471_), .A4(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n476_));
  NOR2_X1   g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(KEYINPUT69), .B2(KEYINPUT8), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n475_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n476_), .B1(new_n475_), .B2(new_n480_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT10), .B(G99gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n465_), .A2(new_n468_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT9), .ZN(new_n487_));
  OAI22_X1  g286(.A1(new_n477_), .A2(KEYINPUT65), .B1(new_n479_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT65), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n489_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n479_), .A2(new_n491_), .A3(new_n487_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n479_), .B2(new_n487_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n488_), .B(new_n490_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT66), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n479_), .A2(new_n487_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT64), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n479_), .A2(new_n491_), .A3(new_n487_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT66), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(new_n488_), .A4(new_n490_), .ZN(new_n501_));
  AOI211_X1 g300(.A(new_n485_), .B(new_n486_), .C1(new_n495_), .C2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n459_), .B1(new_n483_), .B2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n486_), .B1(new_n495_), .B2(new_n501_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n485_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n475_), .A2(new_n480_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n476_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n475_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n506_), .A2(new_n511_), .A3(new_n443_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n503_), .A2(KEYINPUT12), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT12), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n459_), .B(new_n514_), .C1(new_n483_), .C2(new_n502_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n458_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n503_), .A2(new_n512_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n458_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G120gat), .B(G148gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT73), .ZN(new_n522_));
  XOR2_X1   g321(.A(G176gat), .B(G204gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n520_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT74), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n520_), .A2(new_n526_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n520_), .A2(KEYINPUT74), .A3(new_n526_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT13), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G29gat), .B(G36gat), .ZN(new_n534_));
  INV_X1    g333(.A(G43gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(G50gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT83), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n418_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT84), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n539_), .A2(new_n418_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n538_), .B(KEYINPUT15), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n418_), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n541_), .B(KEYINPUT85), .Z(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT84), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n540_), .A2(new_n550_), .A3(new_n542_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n544_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G169gat), .B(G197gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT86), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G113gat), .ZN(new_n555_));
  INV_X1    g354(.A(G141gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n557_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n544_), .A2(new_n549_), .A3(new_n551_), .A4(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n533_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n546_), .B1(new_n502_), .B2(new_n483_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT76), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT75), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT34), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n569_), .A2(KEYINPUT35), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n506_), .A2(new_n511_), .A3(new_n538_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT77), .Z(new_n572_));
  NAND3_X1  g371(.A1(new_n566_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(KEYINPUT35), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n566_), .A2(KEYINPUT35), .A3(new_n569_), .A4(new_n572_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(G134gat), .ZN(new_n579_));
  INV_X1    g378(.A(G162gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n575_), .A2(new_n576_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n581_), .B(KEYINPUT36), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n575_), .A2(new_n586_), .A3(new_n576_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n584_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT37), .B1(new_n589_), .B2(new_n582_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n455_), .A2(new_n563_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n257_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n408_), .A3(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT38), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n589_), .A2(new_n582_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n455_), .A2(new_n563_), .A3(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G1gat), .B1(new_n598_), .B2(new_n257_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(G1324gat));
  OR2_X1    g399(.A1(new_n598_), .A2(new_n336_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(G8gat), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT108), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n336_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n593_), .A2(new_n409_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(KEYINPUT108), .A2(KEYINPUT39), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n601_), .A2(G8gat), .A3(new_n608_), .A4(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n605_), .A2(new_n607_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(G1325gat));
  INV_X1    g412(.A(G15gat), .ZN(new_n614_));
  INV_X1    g413(.A(new_n406_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n593_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G15gat), .B1(new_n598_), .B2(new_n406_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT41), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n616_), .B1(new_n619_), .B2(new_n620_), .ZN(G1326gat));
  INV_X1    g420(.A(G22gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n593_), .A2(new_n622_), .A3(new_n365_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G22gat), .B1(new_n598_), .B2(new_n366_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n624_), .A2(KEYINPUT42), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(KEYINPUT42), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n623_), .B1(new_n625_), .B2(new_n626_), .ZN(G1327gat));
  NOR2_X1   g426(.A1(new_n407_), .A2(new_n597_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n563_), .A2(new_n454_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(G29gat), .B1(new_n631_), .B2(new_n594_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n630_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n405_), .A2(new_n406_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n385_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n637_), .B2(new_n591_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n407_), .A2(KEYINPUT43), .A3(new_n592_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n633_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT44), .B(new_n633_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n642_), .A2(G29gat), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n632_), .B1(new_n644_), .B2(new_n594_), .ZN(G1328gat));
  INV_X1    g444(.A(G36gat), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n628_), .A2(new_n633_), .A3(new_n646_), .A4(new_n606_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT45), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n642_), .A2(new_n606_), .A3(new_n643_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(G36gat), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT109), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT46), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n652_), .A2(new_n653_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n651_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n654_), .A2(new_n657_), .ZN(G1329gat));
  NAND4_X1  g457(.A1(new_n642_), .A2(G43gat), .A3(new_n384_), .A4(new_n643_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n629_), .A2(new_n406_), .A3(new_n630_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(G43gat), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g461(.A1(new_n642_), .A2(new_n365_), .A3(new_n643_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT110), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n664_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(G50gat), .A3(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n631_), .A2(new_n537_), .A3(new_n365_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1331gat));
  INV_X1    g468(.A(KEYINPUT13), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n532_), .B(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n561_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n455_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n597_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n675_), .A2(G57gat), .A3(new_n594_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n673_), .A2(new_n591_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G57gat), .B1(new_n677_), .B2(new_n594_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1332gat));
  INV_X1    g478(.A(G64gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n675_), .B2(new_n606_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT48), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n677_), .A2(new_n680_), .A3(new_n606_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1333gat));
  AOI21_X1  g483(.A(new_n422_), .B1(new_n675_), .B2(new_n615_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT49), .Z(new_n686_));
  NAND3_X1  g485(.A1(new_n677_), .A2(new_n422_), .A3(new_n615_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1334gat));
  NAND3_X1  g487(.A1(new_n677_), .A2(new_n423_), .A3(new_n365_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n423_), .B1(new_n675_), .B2(new_n365_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n691_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(KEYINPUT50), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT50), .B1(new_n692_), .B2(new_n693_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n689_), .B1(new_n694_), .B2(new_n695_), .ZN(G1335gat));
  OR2_X1    g495(.A1(new_n638_), .A2(new_n639_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n672_), .A2(new_n454_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(G85gat), .A3(new_n594_), .ZN(new_n701_));
  INV_X1    g500(.A(G85gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n629_), .A2(new_n698_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n704_), .B2(new_n257_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n701_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(G1336gat));
  AOI21_X1  g507(.A(G92gat), .B1(new_n703_), .B2(new_n606_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n606_), .A2(G92gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n700_), .B2(new_n710_), .ZN(G1337gat));
  OAI211_X1 g510(.A(new_n699_), .B(new_n615_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G99gat), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT114), .ZN(new_n714_));
  INV_X1    g513(.A(new_n384_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(new_n484_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n703_), .A2(new_n716_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n713_), .A2(new_n714_), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n718_), .A2(KEYINPUT113), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(KEYINPUT113), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n713_), .A2(KEYINPUT113), .A3(new_n717_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(G1338gat));
  NAND3_X1  g522(.A1(new_n703_), .A2(new_n353_), .A3(new_n365_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n697_), .A2(new_n365_), .A3(new_n699_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(G106gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(G106gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT53), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT53), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n731_), .B(new_n724_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1339gat));
  NOR2_X1   g532(.A1(new_n606_), .A2(new_n715_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n594_), .A3(new_n366_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT122), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n513_), .A2(new_n458_), .A3(new_n515_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT118), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(KEYINPUT55), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(KEYINPUT55), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n517_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(KEYINPUT55), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT118), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n737_), .A2(new_n738_), .A3(KEYINPUT55), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n516_), .A3(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n741_), .A2(new_n745_), .A3(new_n526_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT119), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT56), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n741_), .A2(new_n745_), .A3(KEYINPUT119), .A4(new_n526_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT120), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n741_), .A2(new_n745_), .A3(KEYINPUT56), .A4(new_n526_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT120), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n748_), .A2(new_n754_), .A3(new_n749_), .A4(new_n750_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n753_), .A3(new_n755_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n561_), .A2(KEYINPUT117), .A3(new_n527_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT117), .B1(new_n561_), .B2(new_n527_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n532_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n540_), .A2(new_n548_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n545_), .A2(new_n547_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n548_), .ZN(new_n764_));
  MUX2_X1   g563(.A(new_n764_), .B(new_n552_), .S(new_n559_), .Z(new_n765_));
  NAND2_X1  g564(.A1(new_n761_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n674_), .B1(new_n760_), .B2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n736_), .B1(new_n767_), .B2(KEYINPUT57), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n756_), .A2(new_n759_), .B1(new_n761_), .B2(new_n765_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NOR4_X1   g569(.A1(new_n769_), .A2(KEYINPUT122), .A3(new_n770_), .A4(new_n674_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n768_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n746_), .A2(new_n749_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n753_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n527_), .A3(new_n765_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT58), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n774_), .A2(new_n765_), .A3(KEYINPUT58), .A4(new_n527_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n591_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT121), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT121), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n777_), .A2(new_n591_), .A3(new_n781_), .A4(new_n778_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n780_), .B(new_n782_), .C1(new_n767_), .C2(KEYINPUT57), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n454_), .B1(new_n772_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n671_), .A2(new_n562_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n454_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n588_), .A2(new_n590_), .A3(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT54), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  OR3_X1    g589(.A1(new_n785_), .A2(new_n787_), .A3(KEYINPUT54), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(KEYINPUT115), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(KEYINPUT115), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n790_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n735_), .B1(new_n784_), .B2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(G113gat), .B1(new_n795_), .B2(new_n561_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n760_), .A2(new_n766_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT57), .A3(new_n597_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT122), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n767_), .A2(new_n736_), .A3(KEYINPUT57), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n783_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n794_), .B1(new_n802_), .B2(new_n786_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n735_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n797_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n735_), .A2(KEYINPUT59), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n779_), .B1(new_n767_), .B2(KEYINPUT57), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n454_), .B1(new_n772_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n809_), .B2(new_n794_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n805_), .A2(new_n562_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n796_), .B1(new_n811_), .B2(G113gat), .ZN(G1340gat));
  XOR2_X1   g611(.A(KEYINPUT123), .B(G120gat), .Z(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n671_), .B2(KEYINPUT60), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n814_), .A2(KEYINPUT60), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n803_), .A2(new_n804_), .A3(new_n815_), .A4(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT124), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n795_), .A2(KEYINPUT124), .A3(new_n815_), .A4(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n808_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n794_), .B1(new_n822_), .B2(new_n786_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n806_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n824_), .B(new_n533_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n813_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n821_), .A2(new_n826_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n795_), .B2(new_n786_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n805_), .A2(new_n810_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n786_), .A2(G127gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT125), .Z(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n829_), .B2(new_n831_), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(new_n795_), .B2(new_n674_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n591_), .A2(G134gat), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT126), .Z(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n829_), .B2(new_n835_), .ZN(G1343gat));
  NOR2_X1   g635(.A1(new_n615_), .A2(new_n366_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n257_), .B(new_n838_), .C1(new_n784_), .C2(new_n794_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n839_), .A2(new_n556_), .A3(new_n561_), .A4(new_n336_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n803_), .A2(new_n594_), .A3(new_n336_), .A4(new_n837_), .ZN(new_n841_));
  OAI21_X1  g640(.A(G141gat), .B1(new_n841_), .B2(new_n562_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1344gat));
  INV_X1    g642(.A(G148gat), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n839_), .A2(new_n844_), .A3(new_n533_), .A4(new_n336_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G148gat), .B1(new_n841_), .B2(new_n671_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1345gat));
  XNOR2_X1  g646(.A(KEYINPUT61), .B(G155gat), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n839_), .A2(new_n336_), .A3(new_n786_), .A4(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n848_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n841_), .B2(new_n454_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1346gat));
  NAND4_X1  g651(.A1(new_n839_), .A2(G162gat), .A3(new_n336_), .A4(new_n591_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n580_), .B1(new_n841_), .B2(new_n597_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1347gat));
  NOR3_X1   g654(.A1(new_n406_), .A2(new_n594_), .A3(new_n336_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n562_), .A2(new_n365_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n823_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G169gat), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n823_), .A2(new_n300_), .A3(new_n856_), .A4(new_n857_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n858_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(G1348gat));
  AND4_X1   g663(.A1(G176gat), .A2(new_n803_), .A3(new_n533_), .A4(new_n366_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n823_), .A2(new_n533_), .A3(new_n366_), .A4(new_n856_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n865_), .A2(new_n856_), .B1(new_n301_), .B2(new_n866_), .ZN(G1349gat));
  AND3_X1   g666(.A1(new_n823_), .A2(new_n366_), .A3(new_n856_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n454_), .A2(new_n296_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n803_), .A2(new_n366_), .A3(new_n786_), .A4(new_n856_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n868_), .A2(new_n869_), .B1(new_n870_), .B2(new_n294_), .ZN(G1350gat));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n591_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G190gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n868_), .A2(new_n292_), .A3(new_n674_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1351gat));
  AOI21_X1  g674(.A(new_n838_), .B1(new_n784_), .B2(new_n794_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n336_), .A2(new_n594_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n561_), .A3(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g678(.A1(new_n876_), .A2(new_n533_), .A3(new_n877_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g680(.A1(new_n876_), .A2(new_n786_), .A3(new_n877_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT63), .B(G211gat), .Z(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n882_), .B2(new_n884_), .ZN(G1354gat));
  NAND3_X1  g684(.A1(new_n876_), .A2(new_n674_), .A3(new_n877_), .ZN(new_n886_));
  INV_X1    g685(.A(G218gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n876_), .A2(G218gat), .A3(new_n591_), .A4(new_n877_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1355gat));
endmodule


