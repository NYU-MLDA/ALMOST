//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT76), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT76), .A2(G155gat), .A3(G162gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT77), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n209_), .A2(new_n214_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n215_));
  OR2_X1    g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n211_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT1), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n213_), .A2(new_n215_), .A3(new_n216_), .A4(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT74), .ZN(new_n226_));
  INV_X1    g025(.A(G127gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(G134gat), .ZN(new_n228_));
  INV_X1    g027(.A(G134gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(G127gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n226_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(G127gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(G134gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT74), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n231_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n223_), .B(KEYINPUT3), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n221_), .B(KEYINPUT2), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n225_), .A2(new_n238_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n238_), .B1(new_n225_), .B2(new_n244_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n225_), .A2(new_n244_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n238_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n220_), .A2(new_n224_), .B1(new_n243_), .B2(new_n241_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n238_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(KEYINPUT4), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n248_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT86), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n246_), .B2(new_n258_), .ZN(new_n259_));
  NOR4_X1   g058(.A1(new_n253_), .A2(new_n238_), .A3(KEYINPUT86), .A4(KEYINPUT4), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n255_), .B(new_n256_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n249_), .B1(new_n261_), .B2(KEYINPUT87), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n248_), .B1(new_n247_), .B2(KEYINPUT4), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT86), .B1(new_n252_), .B2(KEYINPUT4), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n246_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n263_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n206_), .B1(new_n262_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n261_), .A2(KEYINPUT87), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n264_), .A2(new_n267_), .A3(new_n263_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n205_), .A4(new_n249_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT90), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT90), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n275_), .A3(new_n272_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G226gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT19), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT20), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G197gat), .A2(G204gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G197gat), .A2(G204gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT21), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT21), .ZN(new_n291_));
  AND2_X1   g090(.A1(G197gat), .A2(G204gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(new_n287_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294_));
  AND4_X1   g093(.A1(new_n286_), .A2(new_n290_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT80), .B1(new_n290_), .B2(new_n294_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n290_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n295_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(G169gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n301_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT26), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT26), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G190gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT82), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n308_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT25), .B(G183gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n312_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT24), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(G169gat), .B2(G176gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT73), .B1(G169gat), .B2(G176gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320_));
  INV_X1    g119(.A(G169gat), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(new_n319_), .A3(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n302_), .B(KEYINPUT23), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n317_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n306_), .B1(new_n316_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n285_), .B1(new_n299_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n323_), .A2(new_n319_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n317_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n313_), .A2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n331_), .A2(new_n333_), .A3(new_n324_), .A4(new_n325_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n334_), .A2(new_n306_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n290_), .A2(new_n293_), .A3(new_n286_), .A4(new_n294_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n298_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n296_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT83), .B1(new_n335_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT83), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n306_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n299_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n329_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n283_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n284_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n299_), .A2(new_n328_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n344_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n281_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n339_), .A2(new_n342_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n329_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n281_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT20), .B1(new_n299_), .B2(new_n341_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n312_), .A2(new_n315_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n313_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n325_), .B1(G183gat), .B2(G190gat), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n355_), .A2(new_n356_), .B1(new_n357_), .B2(new_n301_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(new_n338_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n283_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n351_), .A2(new_n352_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT85), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n348_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n351_), .A2(new_n360_), .A3(KEYINPUT85), .A4(new_n352_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n338_), .B1(new_n250_), .B2(KEYINPUT29), .ZN(new_n367_));
  XOR2_X1   g166(.A(G22gat), .B(G50gat), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n367_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n253_), .A2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT78), .B(KEYINPUT28), .Z(new_n373_));
  OR2_X1    g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G78gat), .B(G106gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT81), .ZN(new_n376_));
  INV_X1    g175(.A(G233gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n378_), .A2(G228gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(G228gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n377_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n376_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n372_), .A2(new_n373_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n374_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n374_), .B2(new_n384_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n370_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n374_), .A2(new_n384_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n382_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n367_), .B(new_n368_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n374_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT91), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n361_), .A2(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n358_), .B2(new_n338_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n344_), .B1(new_n349_), .B2(new_n397_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n353_), .A2(new_n359_), .A3(new_n283_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n281_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n351_), .A2(new_n360_), .A3(KEYINPUT91), .A4(new_n352_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n395_), .A2(new_n400_), .A3(KEYINPUT27), .A4(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n366_), .A2(new_n393_), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n274_), .A2(new_n276_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT92), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n274_), .A2(new_n403_), .A3(KEYINPUT92), .A4(new_n276_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n393_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n363_), .A2(new_n365_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n267_), .A2(new_n248_), .A3(new_n255_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n205_), .B1(new_n247_), .B2(new_n256_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n262_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT33), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n205_), .A4(new_n270_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n272_), .A2(KEYINPUT33), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n413_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n351_), .A2(new_n360_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n352_), .A2(KEYINPUT32), .ZN(new_n420_));
  OR3_X1    g219(.A1(new_n419_), .A2(KEYINPUT88), .A3(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT88), .B1(new_n419_), .B2(new_n420_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n408_), .B1(new_n418_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n406_), .A2(new_n407_), .A3(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G71gat), .B(G99gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G43gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n341_), .B(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(new_n251_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G227gat), .A2(G233gat), .ZN(new_n432_));
  INV_X1    g231(.A(G15gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT30), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT31), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n431_), .B(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n437_), .B(KEYINPUT75), .Z(new_n438_));
  NAND3_X1  g237(.A1(new_n427_), .A2(KEYINPUT93), .A3(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n274_), .A2(new_n276_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n366_), .A2(new_n402_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n441_), .A2(new_n437_), .A3(new_n393_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT93), .B1(new_n427_), .B2(new_n438_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT71), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT69), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT66), .B(G15gat), .ZN(new_n451_));
  INV_X1    g250(.A(G22gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT67), .B(G8gat), .ZN(new_n454_));
  INV_X1    g253(.A(G1gat), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT14), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT68), .B1(new_n453_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n451_), .B(G22gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n456_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G1gat), .B(G8gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G29gat), .B(G36gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n462_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n464_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n458_), .A2(new_n461_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n462_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n467_), .B1(new_n473_), .B2(new_n463_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n448_), .B(new_n450_), .C1(new_n470_), .C2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n463_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n467_), .B(KEYINPUT15), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n473_), .A2(new_n467_), .A3(new_n463_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n449_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n475_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n468_), .B1(new_n464_), .B2(new_n469_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n479_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n448_), .B1(new_n483_), .B2(new_n450_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G113gat), .B(G141gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT70), .ZN(new_n487_));
  XOR2_X1   g286(.A(G169gat), .B(G197gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n447_), .B1(new_n485_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n450_), .B1(new_n470_), .B2(new_n474_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT69), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n492_), .A2(new_n480_), .A3(new_n475_), .A4(new_n489_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(KEYINPUT71), .ZN(new_n494_));
  OAI22_X1  g293(.A1(new_n490_), .A2(new_n494_), .B1(new_n485_), .B2(new_n489_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT72), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n446_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G230gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G85gat), .B(G92gat), .Z(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT10), .B(G99gat), .Z(new_n501_));
  INV_X1    g300(.A(G106gat), .ZN(new_n502_));
  AOI22_X1  g301(.A1(KEYINPUT9), .A2(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT6), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n503_), .B(new_n505_), .C1(KEYINPUT9), .C2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT7), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n505_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT8), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n500_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n510_), .B2(new_n500_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n507_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n517_));
  XOR2_X1   g316(.A(G71gat), .B(G78gat), .Z(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n517_), .A2(new_n518_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n514_), .A2(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n507_), .B(new_n521_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(KEYINPUT12), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT12), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n514_), .A2(new_n522_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n499_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n498_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G120gat), .B(G148gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT5), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G176gat), .B(G204gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  OR2_X1    g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n534_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT13), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G232gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT34), .ZN(new_n542_));
  OAI22_X1  g341(.A1(new_n514_), .A2(new_n468_), .B1(KEYINPUT35), .B2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n514_), .A2(new_n477_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(KEYINPUT35), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G190gat), .B(G218gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT64), .ZN(new_n550_));
  XOR2_X1   g349(.A(G134gat), .B(G162gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(KEYINPUT36), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n543_), .A2(new_n544_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n546_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n548_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n554_), .B1(new_n548_), .B2(new_n556_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(KEYINPUT36), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n557_), .B2(KEYINPUT65), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n561_), .A3(new_n564_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n521_), .B(new_n569_), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n476_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  XOR2_X1   g372(.A(G127gat), .B(G155gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT16), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n572_), .A2(new_n573_), .A3(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(KEYINPUT17), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n572_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n540_), .A2(new_n568_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n497_), .A2(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n583_), .A2(G1gat), .A3(new_n440_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n584_), .A2(KEYINPUT38), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n446_), .A2(new_n562_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n440_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n495_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n540_), .A2(new_n581_), .A3(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n586_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n584_), .B1(G1gat), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n585_), .B1(new_n591_), .B2(new_n592_), .ZN(G1324gat));
  INV_X1    g392(.A(new_n583_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n441_), .A3(new_n454_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n586_), .A2(new_n589_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n441_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G8gat), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT94), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT94), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n601_), .B(G8gat), .C1(new_n596_), .C2(new_n597_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n599_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n600_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n595_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(G1325gat));
  OAI21_X1  g406(.A(G15gat), .B1(new_n596_), .B2(new_n438_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT41), .Z(new_n609_));
  INV_X1    g408(.A(new_n438_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n594_), .A2(new_n433_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(G1326gat));
  OAI21_X1  g411(.A(G22gat), .B1(new_n596_), .B2(new_n408_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT42), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n594_), .A2(new_n452_), .A3(new_n393_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT95), .Z(G1327gat));
  INV_X1    g416(.A(new_n562_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n581_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n540_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n497_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(G29gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n587_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n539_), .A2(new_n581_), .A3(new_n495_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT43), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n627_), .B(new_n568_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n427_), .A2(new_n438_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT93), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n443_), .A3(new_n439_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n627_), .B1(new_n633_), .B2(new_n568_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n626_), .B1(new_n629_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT44), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n587_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(KEYINPUT96), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n566_), .A2(new_n567_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT43), .B1(new_n446_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n628_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n626_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(KEYINPUT97), .B(KEYINPUT44), .Z(new_n645_));
  AOI21_X1  g444(.A(new_n637_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n623_), .B1(new_n646_), .B2(KEYINPUT98), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n648_));
  INV_X1    g447(.A(new_n645_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n638_), .B2(new_n643_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n648_), .B1(new_n650_), .B2(new_n637_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT99), .B1(new_n647_), .B2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n642_), .B1(new_n641_), .B2(new_n626_), .ZN(new_n653_));
  AOI211_X1 g452(.A(KEYINPUT96), .B(new_n625_), .C1(new_n640_), .C2(new_n628_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n645_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n637_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(KEYINPUT98), .A3(new_n656_), .ZN(new_n657_));
  AND4_X1   g456(.A1(KEYINPUT99), .A2(new_n651_), .A3(new_n657_), .A4(G29gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n624_), .B1(new_n652_), .B2(new_n658_), .ZN(G1328gat));
  INV_X1    g458(.A(G36gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n622_), .A2(new_n660_), .A3(new_n441_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT45), .Z(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n635_), .A2(new_n636_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n650_), .A2(new_n597_), .A3(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n663_), .B(KEYINPUT46), .C1(new_n660_), .C2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT46), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n664_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n660_), .B1(new_n668_), .B2(new_n441_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n669_), .B2(new_n662_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n666_), .A2(new_n670_), .ZN(G1329gat));
  INV_X1    g470(.A(new_n437_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n668_), .A2(G43gat), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G43gat), .B1(new_n622_), .B2(new_n610_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT100), .Z(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT47), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n673_), .A2(new_n675_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1330gat));
  AOI21_X1  g479(.A(G50gat), .B1(new_n622_), .B2(new_n393_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n393_), .A2(G50gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n668_), .B2(new_n682_), .ZN(G1331gat));
  NAND4_X1  g482(.A1(new_n586_), .A2(new_n619_), .A3(new_n540_), .A4(new_n496_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n440_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n446_), .A2(new_n495_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n686_), .A2(new_n619_), .A3(new_n540_), .A4(new_n639_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n440_), .A2(G57gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n685_), .B1(new_n687_), .B2(new_n688_), .ZN(G1332gat));
  OAI21_X1  g488(.A(G64gat), .B1(new_n684_), .B2(new_n597_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT48), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n597_), .A2(G64gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n687_), .B2(new_n692_), .ZN(G1333gat));
  OAI21_X1  g492(.A(G71gat), .B1(new_n684_), .B2(new_n438_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT101), .B(KEYINPUT49), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n438_), .A2(G71gat), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT102), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n687_), .B2(new_n698_), .ZN(G1334gat));
  OAI21_X1  g498(.A(G78gat), .B1(new_n684_), .B2(new_n408_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT50), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n408_), .A2(G78gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n687_), .B2(new_n702_), .ZN(G1335gat));
  NAND2_X1  g502(.A1(new_n540_), .A2(new_n581_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(new_n618_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n686_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G85gat), .B1(new_n707_), .B2(new_n587_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n704_), .A2(new_n495_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n641_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n641_), .B2(new_n710_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n587_), .A2(G85gat), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT104), .Z(new_n715_));
  AOI21_X1  g514(.A(new_n708_), .B1(new_n713_), .B2(new_n715_), .ZN(G1336gat));
  NOR3_X1   g515(.A1(new_n711_), .A2(new_n712_), .A3(new_n597_), .ZN(new_n717_));
  INV_X1    g516(.A(G92gat), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n441_), .A2(new_n718_), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n717_), .A2(new_n718_), .B1(new_n706_), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT105), .ZN(G1337gat));
  AND3_X1   g520(.A1(new_n707_), .A2(new_n501_), .A3(new_n672_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n641_), .A2(new_n710_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n610_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(G99gat), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g525(.A(new_n502_), .B1(new_n723_), .B2(new_n393_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n727_), .A2(KEYINPUT52), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(KEYINPUT52), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n707_), .A2(new_n502_), .A3(new_n393_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT106), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n729_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT53), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n728_), .A2(new_n734_), .A3(new_n729_), .A4(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1339gat));
  INV_X1    g535(.A(G113gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT54), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT108), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n539_), .B(new_n639_), .C1(KEYINPUT108), .C2(new_n738_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n496_), .A2(new_n619_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(KEYINPUT107), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n496_), .A2(new_n744_), .A3(new_n619_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n740_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n742_), .A2(KEYINPUT107), .ZN(new_n747_));
  INV_X1    g546(.A(new_n741_), .ZN(new_n748_));
  AND4_X1   g547(.A1(new_n740_), .A2(new_n747_), .A3(new_n745_), .A4(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n746_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n537_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n485_), .A2(new_n447_), .A3(new_n489_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n493_), .A2(KEYINPUT71), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n489_), .B1(new_n483_), .B2(new_n449_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n478_), .A2(new_n479_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n450_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n756_), .A2(new_n757_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n751_), .A2(new_n754_), .A3(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n525_), .A2(new_n499_), .A3(new_n527_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT55), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(new_n528_), .ZN(new_n765_));
  AOI211_X1 g564(.A(KEYINPUT55), .B(new_n499_), .C1(new_n525_), .C2(new_n527_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n765_), .A2(KEYINPUT110), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n525_), .A2(new_n527_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n498_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(KEYINPUT55), .A3(new_n763_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n766_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n534_), .B1(new_n767_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT110), .B1(new_n765_), .B2(new_n766_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n771_), .A2(new_n772_), .A3(new_n768_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n534_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n776_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n495_), .A2(KEYINPUT109), .A3(new_n535_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT109), .B1(new_n495_), .B2(new_n535_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n762_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(KEYINPUT57), .A3(new_n618_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT57), .B1(new_n785_), .B2(new_n618_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n754_), .A2(new_n535_), .A3(new_n761_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(KEYINPUT112), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n754_), .A2(new_n793_), .A3(new_n535_), .A4(new_n761_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n534_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n534_), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n775_), .B(new_n796_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n794_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n790_), .B1(new_n792_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n791_), .A2(KEYINPUT112), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n781_), .A2(new_n801_), .A3(KEYINPUT113), .A4(new_n794_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(KEYINPUT114), .A3(new_n568_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n781_), .A2(new_n801_), .A3(new_n794_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(new_n800_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT58), .B1(new_n805_), .B2(new_n790_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n639_), .B1(new_n809_), .B2(new_n802_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(KEYINPUT114), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n789_), .B1(new_n808_), .B2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n750_), .B1(new_n812_), .B2(new_n581_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n440_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n442_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n737_), .B1(new_n815_), .B2(new_n588_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT115), .B(new_n737_), .C1(new_n815_), .C2(new_n588_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n814_), .A2(KEYINPUT59), .A3(new_n442_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT116), .B(G113gat), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n496_), .A2(new_n824_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n818_), .A2(new_n819_), .B1(new_n823_), .B2(new_n825_), .ZN(G1340gat));
  AOI21_X1  g625(.A(new_n539_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n827_));
  INV_X1    g626(.A(G120gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n539_), .B2(KEYINPUT60), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(KEYINPUT60), .B2(new_n828_), .ZN(new_n830_));
  OAI22_X1  g629(.A1(new_n827_), .A2(new_n828_), .B1(new_n815_), .B2(new_n830_), .ZN(G1341gat));
  OAI21_X1  g630(.A(new_n227_), .B1(new_n815_), .B2(new_n581_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT117), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n227_), .C1(new_n815_), .C2(new_n581_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n581_), .A2(new_n227_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n833_), .A2(new_n835_), .B1(new_n823_), .B2(new_n836_), .ZN(G1342gat));
  AOI21_X1  g636(.A(new_n639_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n562_), .A2(new_n229_), .ZN(new_n839_));
  OAI22_X1  g638(.A1(new_n838_), .A2(new_n229_), .B1(new_n815_), .B2(new_n839_), .ZN(G1343gat));
  AND2_X1   g639(.A1(new_n438_), .A2(new_n403_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n814_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n495_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g644(.A1(new_n842_), .A2(new_n539_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT118), .B(G148gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1345gat));
  OAI21_X1  g647(.A(KEYINPUT119), .B1(new_n842_), .B2(new_n581_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n814_), .A2(new_n850_), .A3(new_n619_), .A4(new_n841_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n849_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1346gat));
  OR3_X1    g654(.A1(new_n842_), .A2(G162gat), .A3(new_n618_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G162gat), .B1(new_n842_), .B2(new_n639_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1347gat));
  NOR3_X1   g657(.A1(new_n587_), .A2(new_n438_), .A3(new_n393_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n813_), .A2(new_n597_), .A3(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT22), .B(G169gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n495_), .A2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT121), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n861_), .A2(new_n864_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n746_), .A2(new_n749_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n785_), .A2(new_n618_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n786_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n806_), .B1(new_n810_), .B2(KEYINPUT114), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n803_), .A2(new_n568_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n870_), .B1(new_n871_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n866_), .B1(new_n875_), .B2(new_n619_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n876_), .A2(new_n441_), .A3(new_n495_), .A4(new_n859_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n878_), .A3(G169gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n877_), .B2(G169gat), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n880_), .A2(new_n881_), .A3(KEYINPUT62), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n877_), .A2(G169gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT120), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n885_), .B2(new_n879_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n865_), .B1(new_n882_), .B2(new_n886_), .ZN(G1348gat));
  NAND2_X1  g686(.A1(new_n861_), .A2(new_n540_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g688(.A1(new_n861_), .A2(new_n619_), .ZN(new_n890_));
  MUX2_X1   g689(.A(new_n313_), .B(G183gat), .S(new_n890_), .Z(G1350gat));
  NAND2_X1  g690(.A1(new_n861_), .A2(new_n568_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G190gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n861_), .A2(new_n562_), .A3(new_n354_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT122), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n893_), .A2(new_n897_), .A3(new_n894_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1351gat));
  NOR2_X1   g698(.A1(new_n813_), .A2(new_n597_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n587_), .A2(new_n610_), .A3(new_n408_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n903_), .B(new_n495_), .C1(KEYINPUT123), .C2(G197gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT123), .B(G197gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n902_), .B2(new_n588_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1352gat));
  NOR2_X1   g706(.A1(new_n902_), .A2(new_n539_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT124), .B(G204gat), .Z(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1353gat));
  NOR3_X1   g709(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n581_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n912_));
  XOR2_X1   g711(.A(new_n912_), .B(KEYINPUT125), .Z(new_n913_));
  NOR3_X1   g712(.A1(new_n902_), .A2(new_n911_), .A3(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1354gat));
  AND3_X1   g715(.A1(new_n903_), .A2(G218gat), .A3(new_n568_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n902_), .A2(KEYINPUT127), .A3(new_n618_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(G218gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT127), .B1(new_n902_), .B2(new_n618_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n919_), .B2(new_n920_), .ZN(G1355gat));
endmodule


