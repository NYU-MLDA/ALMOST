//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_;
  AND2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT85), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT1), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT86), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n206_), .A2(KEYINPUT1), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(new_n208_), .B2(KEYINPUT86), .ZN(new_n211_));
  AOI211_X1 g010(.A(new_n202_), .B(new_n203_), .C1(new_n209_), .C2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n202_), .A2(KEYINPUT2), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n203_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n202_), .A2(KEYINPUT2), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n213_), .A2(new_n215_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n218_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G113gat), .B(G120gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n221_), .A2(new_n223_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n220_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n212_), .A2(new_n219_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n226_), .A2(KEYINPUT84), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n229_), .B(new_n225_), .Z(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(KEYINPUT98), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT98), .B1(new_n228_), .B2(new_n230_), .ZN(new_n233_));
  OAI211_X1 g032(.A(KEYINPUT4), .B(new_n227_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT99), .B(KEYINPUT4), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n228_), .A2(new_n230_), .A3(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n227_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n233_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(new_n231_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n235_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G1gat), .B(G29gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G85gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT0), .B(G57gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  NAND3_X1  g046(.A1(new_n239_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT100), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n239_), .A2(new_n243_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n239_), .A2(new_n243_), .A3(KEYINPUT100), .A4(new_n247_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G169gat), .ZN(new_n256_));
  INV_X1    g055(.A(G176gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G183gat), .A2(G190gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT23), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(G183gat), .B2(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT94), .ZN(new_n265_));
  OR2_X1    g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n262_), .B1(KEYINPUT24), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n266_), .A2(KEYINPUT24), .A3(new_n259_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT25), .B(G183gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n267_), .A2(new_n268_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n269_), .A2(new_n271_), .A3(new_n274_), .A4(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n265_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G197gat), .B(G204gat), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT21), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT88), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G211gat), .B(G218gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n278_), .B2(KEYINPUT21), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT89), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n283_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n281_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(KEYINPUT21), .A3(new_n286_), .ZN(new_n287_));
  OAI22_X1  g086(.A1(new_n280_), .A2(new_n282_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n277_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n260_), .A2(KEYINPUT82), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n258_), .A2(new_n259_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT82), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n263_), .A3(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n267_), .A2(new_n270_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n274_), .B(KEYINPUT81), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT20), .B1(new_n297_), .B2(new_n288_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n289_), .B1(new_n298_), .B2(KEYINPUT92), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(KEYINPUT92), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G226gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT19), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n299_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n302_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n288_), .B(KEYINPUT91), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(new_n276_), .A3(new_n264_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT20), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n297_), .B2(new_n288_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n304_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n308_), .B(new_n304_), .C1(new_n288_), .C2(new_n277_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT95), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n302_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G64gat), .B(G92gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT97), .ZN(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT96), .B(KEYINPUT18), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G8gat), .B(G36gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT32), .ZN(new_n322_));
  MUX2_X1   g121(.A(new_n310_), .B(new_n314_), .S(new_n322_), .Z(new_n323_));
  NAND2_X1  g122(.A1(new_n255_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT33), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n248_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n314_), .A2(new_n320_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n321_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n248_), .A2(new_n325_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n247_), .B1(new_n242_), .B2(new_n236_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n234_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n326_), .A2(new_n329_), .A3(new_n330_), .A4(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n324_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G22gat), .B(G50gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(G228gat), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n341_));
  NAND2_X1  g140(.A1(new_n228_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n305_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n340_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n288_), .B(new_n340_), .C1(new_n220_), .C2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n336_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n220_), .A2(new_n349_), .A3(new_n345_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n349_), .B1(new_n220_), .B2(new_n345_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353_));
  OR3_X1    g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n336_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n341_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n220_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(new_n305_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n346_), .B(new_n355_), .C1(new_n358_), .C2(new_n340_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n353_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n348_), .A2(new_n354_), .A3(new_n359_), .A4(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n348_), .A2(new_n359_), .B1(new_n354_), .B2(new_n360_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT83), .B(G43gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n297_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(new_n230_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(G15gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT30), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT31), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n369_), .B(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n364_), .A2(new_n375_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n362_), .A2(new_n363_), .A3(new_n375_), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n369_), .B(new_n374_), .Z(new_n378_));
  NAND2_X1  g177(.A1(new_n348_), .A2(new_n359_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n354_), .A2(new_n360_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n378_), .B1(new_n381_), .B2(new_n361_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(new_n255_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n310_), .A2(new_n321_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT27), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n327_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT101), .B1(new_n329_), .B2(KEYINPUT27), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT101), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(new_n386_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n387_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n335_), .A2(new_n376_), .B1(new_n384_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G85gat), .ZN(new_n393_));
  INV_X1    g192(.A(G92gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(G85gat), .A2(G92gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT8), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(G99gat), .A2(G106gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT65), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT7), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT7), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT65), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n400_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  AOI211_X1 g204(.A(G99gat), .B(G106gat), .C1(new_n401_), .C2(KEYINPUT7), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n408_), .B1(G99gat), .B2(G106gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G99gat), .A2(G106gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(KEYINPUT6), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n399_), .B1(new_n407_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n397_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT66), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n410_), .A2(KEYINPUT6), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n408_), .A2(G99gat), .A3(G106gat), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n420_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n418_), .A2(new_n419_), .A3(new_n417_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n416_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n415_), .B1(new_n423_), .B2(new_n398_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT9), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n412_), .B1(new_n425_), .B2(new_n395_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n397_), .A2(KEYINPUT9), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT64), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT10), .B(G99gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(G106gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n429_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n426_), .B(new_n427_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G29gat), .B(G36gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G43gat), .B(G50gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n424_), .A2(new_n434_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT66), .B1(new_n409_), .B2(new_n411_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n400_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n403_), .A2(KEYINPUT65), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n401_), .A2(KEYINPUT7), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n402_), .A2(new_n400_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n439_), .A2(new_n422_), .A3(new_n443_), .A4(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n398_), .B1(new_n445_), .B2(new_n397_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n434_), .B1(new_n446_), .B2(new_n414_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n437_), .B(KEYINPUT15), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT73), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G232gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT34), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT35), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n450_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n438_), .A2(new_n449_), .A3(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n453_), .A2(new_n454_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n457_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n438_), .A2(new_n449_), .A3(new_n459_), .A4(new_n455_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G190gat), .B(G218gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(G134gat), .B(G162gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(KEYINPUT36), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n461_), .A2(KEYINPUT72), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n458_), .A2(KEYINPUT72), .A3(new_n460_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(KEYINPUT36), .B2(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n467_), .A2(KEYINPUT36), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n461_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n392_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G8gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT74), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G1gat), .A2(G8gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT14), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n478_), .A2(KEYINPUT74), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n478_), .A2(KEYINPUT74), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n482_), .A3(new_n480_), .A4(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G231gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT67), .B(G71gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G78gat), .ZN(new_n492_));
  OR2_X1    g291(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n493_));
  INV_X1    g292(.A(G78gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n492_), .A2(new_n496_), .B1(KEYINPUT11), .B2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(KEYINPUT11), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n492_), .A2(new_n496_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n490_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT75), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT76), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT76), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n503_), .A2(new_n504_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G127gat), .B(G155gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT16), .ZN(new_n511_));
  XOR2_X1   g310(.A(G183gat), .B(G211gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(KEYINPUT17), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT17), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n503_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n516_), .B2(new_n513_), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n509_), .B(new_n517_), .Z(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G230gat), .A2(G233gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n447_), .A2(new_n502_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n434_), .B(new_n501_), .C1(new_n446_), .C2(new_n414_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT12), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n521_), .A2(new_n522_), .B1(new_n524_), .B2(new_n447_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT69), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n501_), .B1(new_n424_), .B2(new_n434_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n521_), .A2(KEYINPUT69), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n525_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n523_), .B1(new_n532_), .B2(new_n520_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G120gat), .B(G148gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT5), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n533_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT13), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n488_), .A2(new_n437_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n437_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n484_), .A2(new_n545_), .A3(new_n487_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT77), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n437_), .B(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n544_), .B(new_n543_), .C1(new_n550_), .C2(new_n488_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT78), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n448_), .A2(new_n487_), .A3(new_n484_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT78), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(new_n544_), .A3(new_n554_), .A4(new_n543_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n548_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G169gat), .B(G197gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n548_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n562_), .A2(KEYINPUT79), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT79), .B1(new_n562_), .B2(new_n563_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n542_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n477_), .A2(new_n519_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n255_), .ZN(new_n571_));
  OAI21_X1  g370(.A(G1gat), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT103), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT103), .B(G1gat), .C1(new_n570_), .C2(new_n571_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT80), .ZN(new_n577_));
  INV_X1    g376(.A(new_n565_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n562_), .A2(KEYINPUT79), .A3(new_n563_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n564_), .A2(new_n565_), .A3(KEYINPUT80), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n474_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(new_n518_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n542_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n377_), .A2(new_n382_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n391_), .A2(new_n590_), .A3(new_n571_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n376_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n324_), .B2(new_n334_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n582_), .B(new_n589_), .C1(new_n591_), .C2(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT102), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(KEYINPUT102), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n571_), .A2(G1gat), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT38), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n595_), .A2(new_n600_), .A3(new_n596_), .A4(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n576_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT104), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n576_), .A2(new_n602_), .A3(KEYINPUT104), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(G1324gat));
  NAND2_X1  g406(.A1(new_n595_), .A2(new_n596_), .ZN(new_n608_));
  OR3_X1    g407(.A1(new_n608_), .A2(G8gat), .A3(new_n391_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G8gat), .B1(new_n570_), .B2(new_n391_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(KEYINPUT39), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(KEYINPUT39), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n609_), .B(new_n614_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1325gat));
  OAI21_X1  g417(.A(G15gat), .B1(new_n570_), .B2(new_n378_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n620_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n375_), .A2(new_n371_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n621_), .B(new_n622_), .C1(new_n608_), .C2(new_n623_), .ZN(G1326gat));
  INV_X1    g423(.A(new_n364_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G22gat), .B1(new_n570_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT42), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n625_), .A2(G22gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n627_), .B1(new_n608_), .B2(new_n628_), .ZN(G1327gat));
  INV_X1    g428(.A(KEYINPUT43), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n583_), .B(KEYINPUT37), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n630_), .B1(new_n392_), .B2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(KEYINPUT43), .B(new_n585_), .C1(new_n591_), .C2(new_n593_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n632_), .A2(new_n518_), .A3(new_n633_), .A4(new_n569_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n585_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n519_), .B1(new_n637_), .B2(new_n630_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n638_), .A2(KEYINPUT44), .A3(new_n569_), .A4(new_n633_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n636_), .A2(new_n639_), .A3(G29gat), .A4(new_n255_), .ZN(new_n640_));
  INV_X1    g439(.A(G29gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n582_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n392_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n518_), .A2(new_n476_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n588_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n641_), .B1(new_n646_), .B2(new_n571_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n640_), .A2(new_n647_), .ZN(G1328gat));
  INV_X1    g447(.A(new_n391_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n636_), .A2(new_n639_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G36gat), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n391_), .A2(G36gat), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n646_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT45), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n651_), .A2(new_n655_), .A3(KEYINPUT46), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1329gat));
  INV_X1    g459(.A(G43gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(new_n646_), .B2(new_n378_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n636_), .A2(new_n639_), .A3(G43gat), .A4(new_n375_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT47), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT47), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(new_n668_), .A3(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1330gat));
  OR3_X1    g469(.A1(new_n646_), .A2(G50gat), .A3(new_n625_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n636_), .A2(new_n639_), .A3(new_n364_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n672_), .A2(new_n673_), .A3(G50gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n672_), .B2(G50gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(G1331gat));
  NOR3_X1   g475(.A1(new_n542_), .A2(new_n582_), .A3(new_n518_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n477_), .A2(new_n255_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G57gat), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n392_), .A2(new_n567_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(new_n588_), .A3(new_n586_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n571_), .A2(G57gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(G1332gat));
  OR3_X1    g482(.A1(new_n681_), .A2(G64gat), .A3(new_n391_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n477_), .A2(new_n649_), .A3(new_n677_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G64gat), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(KEYINPUT48), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(KEYINPUT48), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1333gat));
  OR3_X1    g488(.A1(new_n681_), .A2(G71gat), .A3(new_n378_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n477_), .A2(new_n375_), .A3(new_n677_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G71gat), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(KEYINPUT49), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(KEYINPUT49), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(G1334gat));
  NAND3_X1  g494(.A1(new_n477_), .A2(new_n364_), .A3(new_n677_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G78gat), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT50), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT50), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n364_), .A2(new_n494_), .ZN(new_n700_));
  OAI22_X1  g499(.A1(new_n698_), .A2(new_n699_), .B1(new_n681_), .B2(new_n700_), .ZN(G1335gat));
  NOR2_X1   g500(.A1(new_n542_), .A2(new_n567_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n632_), .A2(new_n518_), .A3(new_n633_), .A4(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n571_), .ZN(new_n704_));
  NOR4_X1   g503(.A1(new_n392_), .A2(new_n567_), .A3(new_n542_), .A4(new_n644_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n393_), .A3(new_n255_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1336gat));
  OAI21_X1  g506(.A(G92gat), .B1(new_n703_), .B2(new_n391_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n705_), .A2(new_n394_), .A3(new_n649_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1337gat));
  OAI21_X1  g509(.A(G99gat), .B1(new_n703_), .B2(new_n378_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n705_), .A2(new_n430_), .A3(new_n375_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g513(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n715_));
  OAI21_X1  g514(.A(G106gat), .B1(new_n703_), .B2(new_n625_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT52), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n718_), .B(G106gat), .C1(new_n703_), .C2(new_n625_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n625_), .A2(G106gat), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n705_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n715_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n722_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n715_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n724_), .B(new_n725_), .C1(new_n717_), .C2(new_n719_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1339gat));
  INV_X1    g526(.A(new_n540_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT111), .B1(new_n532_), .B2(new_n520_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n447_), .A2(new_n524_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n522_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n527_), .B2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT69), .B1(new_n521_), .B2(new_n530_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n526_), .B(new_n528_), .C1(new_n447_), .C2(new_n502_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n736_), .A2(new_n737_), .A3(G230gat), .A4(G233gat), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n529_), .A2(new_n531_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n739_), .A2(KEYINPUT55), .A3(new_n520_), .A4(new_n733_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n733_), .B(new_n520_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n730_), .A2(new_n738_), .A3(new_n740_), .A4(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n537_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n537_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n729_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n544_), .A2(new_n546_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n560_), .B1(new_n749_), .B2(new_n543_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n553_), .A2(new_n544_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n543_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n563_), .A2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(KEYINPUT112), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n563_), .B2(new_n752_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n541_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n476_), .B1(new_n748_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT57), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n540_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n744_), .A2(new_n537_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT56), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n764_), .B2(new_n745_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n757_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n583_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n540_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n764_), .B2(new_n745_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n631_), .B1(new_n769_), .B2(KEYINPUT58), .ZN(new_n770_));
  INV_X1    g569(.A(new_n768_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n760_), .A2(new_n767_), .B1(new_n770_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n759_), .B1(new_n775_), .B2(KEYINPUT115), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n771_), .B(KEYINPUT58), .C1(new_n746_), .C2(new_n747_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n773_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n777_), .B(new_n585_), .C1(new_n769_), .C2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(KEYINPUT115), .C1(KEYINPUT57), .C2(new_n758_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n518_), .B1(new_n776_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n586_), .A2(new_n642_), .A3(new_n542_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT54), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n391_), .A2(new_n255_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n786_), .A2(new_n378_), .A3(new_n364_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n519_), .B1(new_n775_), .B2(new_n759_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n783_), .B(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n779_), .B1(KEYINPUT57), .B2(new_n758_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n767_), .A2(new_n760_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n518_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n784_), .A3(KEYINPUT114), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n795_), .A2(new_n799_), .A3(new_n787_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n790_), .B1(new_n800_), .B2(new_n788_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G113gat), .B1(new_n801_), .B2(new_n642_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n795_), .A2(new_n799_), .A3(new_n787_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n804_), .A2(G113gat), .A3(new_n566_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n802_), .A2(new_n803_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(G113gat), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n804_), .A2(KEYINPUT59), .B1(new_n785_), .B2(new_n789_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n582_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT116), .B1(new_n810_), .B2(new_n805_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n807_), .A2(new_n811_), .ZN(G1340gat));
  OAI21_X1  g611(.A(G120gat), .B1(new_n801_), .B2(new_n542_), .ZN(new_n813_));
  INV_X1    g612(.A(G120gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n542_), .B2(KEYINPUT60), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(KEYINPUT60), .B2(new_n814_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n813_), .B1(new_n804_), .B2(new_n816_), .ZN(G1341gat));
  AOI21_X1  g616(.A(G127gat), .B1(new_n800_), .B2(new_n519_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n519_), .A2(G127gat), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n819_), .B(KEYINPUT117), .Z(new_n820_));
  AOI21_X1  g619(.A(new_n818_), .B1(new_n809_), .B2(new_n820_), .ZN(G1342gat));
  AOI21_X1  g620(.A(G134gat), .B1(new_n800_), .B2(new_n476_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n585_), .A2(G134gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT118), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n809_), .B2(new_n824_), .ZN(G1343gat));
  NAND2_X1  g624(.A1(new_n795_), .A2(new_n799_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n826_), .A2(new_n375_), .A3(new_n625_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n786_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT119), .B(G141gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n567_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n831_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n829_), .B2(new_n566_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1344gat));
  OR3_X1    g634(.A1(new_n829_), .A2(G148gat), .A3(new_n542_), .ZN(new_n836_));
  OAI21_X1  g635(.A(G148gat), .B1(new_n829_), .B2(new_n542_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1345gat));
  XNOR2_X1  g637(.A(KEYINPUT61), .B(G155gat), .ZN(new_n839_));
  OR3_X1    g638(.A1(new_n829_), .A2(new_n518_), .A3(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n829_), .B2(new_n518_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1346gat));
  INV_X1    g641(.A(G162gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n631_), .A2(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT120), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n827_), .A2(new_n476_), .A3(new_n828_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n830_), .A2(new_n845_), .B1(new_n846_), .B2(new_n843_), .ZN(G1347gat));
  NOR2_X1   g646(.A1(new_n391_), .A2(new_n255_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n382_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n567_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n852_));
  INV_X1    g651(.A(new_n256_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n851_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT62), .B1(new_n851_), .B2(G169gat), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1348gat));
  NAND2_X1  g655(.A1(new_n848_), .A2(new_n375_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(G176gat), .A3(new_n588_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n795_), .A2(new_n625_), .A3(new_n799_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n795_), .A2(new_n799_), .A3(KEYINPUT121), .A4(new_n625_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n859_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  AOI21_X1  g664(.A(G176gat), .B1(new_n850_), .B2(new_n588_), .ZN(new_n866_));
  OR3_X1    g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1349gat));
  NOR2_X1   g668(.A1(new_n518_), .A2(new_n272_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n850_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n858_), .A2(new_n519_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(G183gat), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(new_n871_), .C1(new_n873_), .C2(G183gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1350gat));
  NAND2_X1  g677(.A1(new_n850_), .A2(new_n585_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(G190gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n850_), .A2(new_n476_), .A3(new_n273_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1351gat));
  INV_X1    g681(.A(new_n826_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n377_), .A3(new_n848_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n885_), .A2(KEYINPUT124), .A3(G197gat), .A4(new_n567_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n883_), .A2(new_n377_), .A3(new_n567_), .A4(new_n848_), .ZN(new_n888_));
  INV_X1    g687(.A(G197gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n889_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n886_), .A2(new_n890_), .A3(new_n891_), .ZN(G1352gat));
  OAI22_X1  g691(.A1(new_n884_), .A2(new_n542_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n893_));
  NAND2_X1  g692(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT126), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n893_), .B(new_n895_), .ZN(G1353gat));
  XOR2_X1   g695(.A(KEYINPUT63), .B(G211gat), .Z(new_n897_));
  NAND3_X1  g696(.A1(new_n885_), .A2(new_n519_), .A3(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n884_), .B2(new_n518_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1354gat));
  AOI21_X1  g700(.A(G218gat), .B1(new_n885_), .B2(new_n476_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n585_), .A2(G218gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT127), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n885_), .B2(new_n904_), .ZN(G1355gat));
endmodule


