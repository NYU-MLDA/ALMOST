//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT9), .ZN(new_n205_));
  NOR3_X1   g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT10), .B(G99gat), .Z(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n203_), .A2(new_n205_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n212_), .A2(KEYINPUT64), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218_));
  AND3_X1   g017(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G92gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT9), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n221_), .A2(new_n226_), .A3(new_n216_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT10), .B(G99gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(G106gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n218_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n217_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G57gat), .ZN(new_n232_));
  INV_X1    g031(.A(G64gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G57gat), .A2(G64gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n237_));
  INV_X1    g036(.A(G78gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n238_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n242_));
  OAI211_X1 g041(.A(KEYINPUT11), .B(new_n236_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n234_), .A2(new_n246_), .A3(new_n235_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n244_), .A2(new_n245_), .A3(new_n247_), .A4(new_n240_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n203_), .A2(new_n204_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT7), .ZN(new_n251_));
  INV_X1    g050(.A(G99gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(new_n252_), .A3(new_n214_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n250_), .B1(new_n255_), .B2(new_n211_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT8), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n255_), .A2(KEYINPUT65), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n221_), .B1(new_n255_), .B2(KEYINPUT65), .ZN(new_n260_));
  OAI211_X1 g059(.A(KEYINPUT8), .B(new_n250_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n231_), .A2(new_n249_), .A3(new_n258_), .A4(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT12), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n217_), .A2(new_n230_), .B1(new_n257_), .B2(new_n256_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n249_), .B1(new_n264_), .B2(new_n261_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  AOI211_X1 g065(.A(KEYINPUT12), .B(new_n249_), .C1(new_n264_), .C2(new_n261_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n202_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n231_), .A2(new_n258_), .A3(new_n261_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n249_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n262_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n202_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(KEYINPUT67), .A3(new_n271_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n268_), .A2(new_n269_), .A3(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G120gat), .B(G148gat), .ZN(new_n279_));
  INV_X1    g078(.A(G204gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT5), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(G176gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT69), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n274_), .A2(KEYINPUT68), .A3(new_n275_), .A4(new_n276_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n278_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n283_), .B1(new_n278_), .B2(new_n285_), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT70), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n278_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n290_));
  INV_X1    g089(.A(new_n285_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n272_), .A2(KEYINPUT12), .A3(new_n262_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n263_), .A2(new_n265_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n275_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(KEYINPUT68), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n291_), .B1(new_n295_), .B2(new_n277_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n289_), .B(new_n290_), .C1(new_n296_), .C2(new_n283_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n288_), .A2(KEYINPUT13), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT13), .B1(new_n288_), .B2(new_n297_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G78gat), .B(G106gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G228gat), .A2(G233gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT88), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308_));
  AND2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT89), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n308_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT89), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n307_), .B(new_n313_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G141gat), .B(G148gat), .Z(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OR4_X1    g116(.A1(KEYINPUT90), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n322_));
  OAI22_X1  g121(.A1(KEYINPUT90), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n318_), .A2(new_n321_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n309_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n307_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n317_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT29), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G211gat), .B(G218gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT93), .ZN(new_n330_));
  INV_X1    g129(.A(G197gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(G204gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n280_), .A2(G197gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT21), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT92), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n331_), .B2(G204gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n280_), .A2(KEYINPUT92), .A3(G197gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT21), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n330_), .A2(new_n334_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT94), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n342_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n330_), .A2(new_n339_), .A3(new_n338_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n305_), .B1(new_n328_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(new_n317_), .B2(new_n326_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n346_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n305_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n304_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G22gat), .B(G50gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n327_), .B2(KEYINPUT29), .ZN(new_n358_));
  INV_X1    g157(.A(new_n357_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n317_), .A2(new_n350_), .A3(new_n326_), .A4(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n356_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n328_), .A2(new_n305_), .A3(new_n348_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n353_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n304_), .B(KEYINPUT95), .Z(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n358_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n355_), .A2(new_n362_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT96), .ZN(new_n369_));
  INV_X1    g168(.A(new_n366_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n365_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n367_), .ZN(new_n372_));
  OAI22_X1  g171(.A1(new_n370_), .A2(new_n371_), .B1(new_n372_), .B2(new_n361_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n361_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT96), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n366_), .A4(new_n355_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n369_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT23), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT79), .B(G183gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT80), .B(G190gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(G176gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT22), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT83), .B1(new_n390_), .B2(G169gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT22), .B(G169gat), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n389_), .B(new_n391_), .C1(new_n392_), .C2(KEYINPUT83), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n387_), .A2(new_n388_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n385_), .A2(KEYINPUT25), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(KEYINPUT25), .B2(G183gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT26), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G190gat), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n396_), .B(new_n398_), .C1(new_n397_), .C2(new_n386_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(G169gat), .A2(G176gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n400_), .B(KEYINPUT81), .Z(new_n401_));
  OR2_X1    g200(.A1(new_n401_), .A2(KEYINPUT24), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(KEYINPUT24), .A3(new_n388_), .ZN(new_n403_));
  MUX2_X1   g202(.A(new_n378_), .B(new_n380_), .S(new_n382_), .Z(new_n404_));
  NAND4_X1  g203(.A1(new_n399_), .A2(new_n402_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n394_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT87), .B(G127gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G134gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G113gat), .B(G120gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT31), .ZN(new_n411_));
  AND2_X1   g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n412_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n406_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n414_), .A3(new_n406_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G71gat), .B(G99gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT85), .ZN(new_n419_));
  XOR2_X1   g218(.A(KEYINPUT86), .B(KEYINPUT30), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G15gat), .B(G43gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT84), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n421_), .B(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n416_), .A2(new_n417_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n413_), .A2(new_n414_), .A3(new_n406_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n415_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n377_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n428_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n431_), .A2(new_n369_), .A3(new_n373_), .A4(new_n376_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n410_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n327_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n317_), .A2(new_n410_), .A3(new_n326_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G1gat), .B(G29gat), .Z(new_n440_));
  XNOR2_X1  g239(.A(G57gat), .B(G85gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n442_), .B(new_n443_), .Z(new_n444_));
  OR2_X1    g243(.A1(new_n435_), .A2(KEYINPUT4), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n435_), .A2(KEYINPUT4), .A3(new_n436_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n439_), .B(new_n444_), .C1(new_n447_), .C2(new_n438_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n444_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n438_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n439_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G226gat), .A2(G233gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n455_), .B(KEYINPUT97), .Z(new_n456_));
  XOR2_X1   g255(.A(new_n456_), .B(KEYINPUT19), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT20), .B1(new_n348_), .B2(new_n406_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n404_), .B1(G183gat), .B2(G190gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n392_), .A2(new_n389_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n388_), .A3(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT25), .B(G183gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT26), .B(G190gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n388_), .A2(KEYINPUT24), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n466_), .A2(KEYINPUT98), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(KEYINPUT98), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n401_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT24), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n400_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n384_), .A2(new_n465_), .A3(new_n469_), .A4(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n462_), .A2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n352_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n458_), .B1(new_n459_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n473_), .B2(new_n352_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n348_), .A2(new_n406_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n457_), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT18), .B(G64gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(G92gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G8gat), .B(G36gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n479_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT101), .ZN(new_n485_));
  INV_X1    g284(.A(new_n483_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n459_), .A2(new_n474_), .A3(new_n458_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n457_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT101), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n475_), .A2(new_n479_), .A3(new_n490_), .A4(new_n483_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n485_), .A2(KEYINPUT27), .A3(new_n489_), .A4(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT27), .ZN(new_n493_));
  INV_X1    g292(.A(new_n484_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n483_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n433_), .A2(new_n454_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n438_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n437_), .A2(new_n500_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n501_), .B(KEYINPUT33), .C1(new_n447_), .C2(new_n500_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n444_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n494_), .A2(new_n495_), .ZN(new_n504_));
  OAI211_X1 g303(.A(KEYINPUT33), .B(new_n449_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n505_));
  OR3_X1    g304(.A1(new_n450_), .A2(KEYINPUT33), .A3(new_n451_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .A4(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n483_), .A2(KEYINPUT32), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n509_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT100), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n475_), .A2(new_n479_), .A3(new_n508_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT100), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n513_), .B(new_n509_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n453_), .A2(new_n511_), .A3(new_n512_), .A4(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n377_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n429_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n499_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G232gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT34), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT15), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT72), .B(G43gat), .ZN(new_n523_));
  INV_X1    g322(.A(G50gat), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G29gat), .B(G36gat), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n524_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n526_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n522_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n523_), .B(new_n524_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n526_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(KEYINPUT15), .A3(new_n528_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n531_), .A2(new_n535_), .B1(new_n264_), .B2(new_n261_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n528_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n270_), .A2(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(KEYINPUT35), .B(new_n521_), .C1(new_n536_), .C2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n531_), .A2(new_n535_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n270_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n521_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n543_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n264_), .A2(new_n528_), .A3(new_n534_), .A4(new_n261_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n541_), .A2(new_n545_), .A3(new_n546_), .A4(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n539_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT73), .B(G190gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(G218gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(G134gat), .B(G162gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT36), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n550_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n539_), .A2(new_n548_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT36), .A3(new_n554_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n556_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n557_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G15gat), .B(G22gat), .ZN(new_n562_));
  INV_X1    g361(.A(G1gat), .ZN(new_n563_));
  INV_X1    g362(.A(G8gat), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT14), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G1gat), .B(G8gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n249_), .B(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT76), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n576_), .A2(new_n577_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n571_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n580_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n560_), .A2(new_n561_), .A3(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n519_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n540_), .A2(new_n568_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n537_), .A2(new_n568_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT77), .Z(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n537_), .A2(new_n568_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n591_), .B1(new_n594_), .B2(new_n589_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(G113gat), .B(G141gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(G169gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(new_n331_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n593_), .A2(new_n595_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT78), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n600_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n596_), .A2(KEYINPUT78), .A3(new_n599_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n303_), .A2(new_n587_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(new_n563_), .A3(new_n453_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT103), .ZN(new_n613_));
  INV_X1    g412(.A(new_n585_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n556_), .A2(new_n559_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n499_), .B2(new_n518_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n300_), .A2(new_n606_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n563_), .B1(new_n620_), .B2(new_n453_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n610_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(KEYINPUT102), .A3(KEYINPUT38), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n624_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n621_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n613_), .A2(new_n626_), .ZN(G1324gat));
  NAND3_X1  g426(.A1(new_n618_), .A2(new_n619_), .A3(new_n497_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n628_), .A2(new_n629_), .A3(G8gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n628_), .B2(G8gat), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n497_), .A2(new_n564_), .ZN(new_n632_));
  OAI22_X1  g431(.A1(new_n630_), .A2(new_n631_), .B1(new_n608_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT104), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT104), .ZN(new_n635_));
  OAI221_X1 g434(.A(new_n635_), .B1(new_n608_), .B2(new_n632_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g437(.A(G15gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n620_), .B2(new_n431_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT41), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n609_), .A2(new_n639_), .A3(new_n431_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n620_), .B2(new_n377_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT42), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n609_), .A2(new_n644_), .A3(new_n377_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1327gat));
  AOI21_X1  g447(.A(new_n497_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n377_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n649_), .A2(new_n454_), .B1(new_n650_), .B2(new_n429_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n651_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n619_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G29gat), .B1(new_n654_), .B2(new_n453_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n560_), .A2(new_n561_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n519_), .B2(new_n658_), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT43), .B(new_n657_), .C1(new_n499_), .C2(new_n518_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n619_), .B(new_n585_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT43), .B1(new_n651_), .B2(new_n657_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n519_), .A2(new_n656_), .A3(new_n658_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n666_), .A2(KEYINPUT44), .A3(new_n619_), .A4(new_n585_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n663_), .A2(new_n453_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n655_), .B1(new_n668_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g468(.A1(new_n663_), .A2(new_n497_), .A3(new_n667_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G36gat), .ZN(new_n671_));
  INV_X1    g470(.A(G36gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n652_), .A2(new_n672_), .A3(new_n619_), .ZN(new_n673_));
  OR3_X1    g472(.A1(new_n673_), .A2(KEYINPUT45), .A3(new_n498_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT45), .B1(new_n673_), .B2(new_n498_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n671_), .A2(KEYINPUT46), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  NOR3_X1   g480(.A1(new_n653_), .A2(G43gat), .A3(new_n429_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n663_), .A2(new_n431_), .A3(new_n667_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n683_), .B2(G43gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g484(.A1(new_n663_), .A2(new_n377_), .A3(new_n667_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT105), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT105), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(G50gat), .A3(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n654_), .A2(new_n524_), .A3(new_n377_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1331gat));
  INV_X1    g490(.A(new_n300_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n607_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n587_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n453_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT106), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n302_), .A2(new_n606_), .A3(new_n618_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT107), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n302_), .A2(new_n699_), .A3(new_n618_), .A4(new_n606_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n454_), .A2(new_n232_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n696_), .B1(new_n701_), .B2(new_n702_), .ZN(G1332gat));
  NAND3_X1  g502(.A1(new_n694_), .A2(new_n233_), .A3(new_n497_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n497_), .A3(new_n700_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G64gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n705_), .A2(new_n708_), .A3(G64gat), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n707_), .A2(KEYINPUT48), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT48), .B1(new_n707_), .B2(new_n709_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n704_), .B1(new_n710_), .B2(new_n711_), .ZN(G1333gat));
  INV_X1    g511(.A(G71gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n694_), .A2(new_n713_), .A3(new_n431_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT49), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n701_), .A2(new_n431_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(G71gat), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT49), .B(new_n713_), .C1(new_n701_), .C2(new_n431_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1334gat));
  NAND3_X1  g518(.A1(new_n694_), .A2(new_n238_), .A3(new_n377_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n698_), .A2(new_n377_), .A3(new_n700_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(G78gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n721_), .B2(G78gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT109), .B(new_n720_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1335gat));
  NAND2_X1  g528(.A1(new_n693_), .A2(new_n585_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT110), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n693_), .A2(new_n732_), .A3(new_n585_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n666_), .A2(new_n731_), .A3(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(G85gat), .A3(new_n453_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n303_), .A2(new_n607_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n652_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n222_), .B1(new_n737_), .B2(new_n454_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1336gat));
  NAND3_X1  g538(.A1(new_n734_), .A2(G92gat), .A3(new_n497_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n223_), .B1(new_n737_), .B2(new_n498_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1337gat));
  INV_X1    g541(.A(new_n737_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(new_n213_), .A3(new_n431_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n734_), .A2(new_n431_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n252_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT51), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n744_), .C1(new_n745_), .C2(new_n252_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n743_), .A2(new_n214_), .A3(new_n377_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n666_), .A2(new_n377_), .A3(new_n731_), .A4(new_n733_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G106gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G106gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n751_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1339gat));
  OAI211_X1 g559(.A(new_n586_), .B(new_n606_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n592_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n588_), .A2(new_n590_), .A3(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n592_), .B1(new_n594_), .B2(new_n589_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n599_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT112), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n765_), .A2(new_n769_), .A3(new_n599_), .A4(new_n766_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n602_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n288_), .A2(new_n297_), .A3(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n288_), .A2(new_n297_), .A3(KEYINPUT113), .A4(new_n772_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n268_), .B1(KEYINPUT111), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n292_), .A2(new_n293_), .A3(new_n275_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n294_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n284_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT56), .B(new_n284_), .C1(new_n778_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n278_), .A2(new_n285_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n283_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n607_), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n775_), .A2(new_n776_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n616_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT57), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(KEYINPUT57), .A3(new_n616_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n789_), .A2(new_n772_), .A3(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT114), .B1(new_n287_), .B2(new_n771_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n786_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(KEYINPUT58), .A3(new_n786_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n658_), .A3(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n794_), .A2(new_n795_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n763_), .B1(new_n805_), .B2(new_n585_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n497_), .A2(new_n454_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n806_), .A2(new_n432_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G113gat), .B1(new_n809_), .B2(new_n607_), .ZN(new_n810_));
  INV_X1    g609(.A(G113gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n607_), .B2(KEYINPUT115), .ZN(new_n812_));
  INV_X1    g611(.A(new_n763_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n791_), .A2(KEYINPUT57), .A3(new_n616_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT57), .B1(new_n791_), .B2(new_n616_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n802_), .A2(new_n658_), .A3(new_n803_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n814_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n813_), .B1(new_n817_), .B2(new_n614_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n818_), .A2(new_n517_), .A3(new_n431_), .A4(new_n807_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n809_), .A2(KEYINPUT59), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n812_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n811_), .A2(KEYINPUT115), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n810_), .B1(new_n823_), .B2(new_n824_), .ZN(G1340gat));
  INV_X1    g624(.A(G120gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n692_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n809_), .B(new_n827_), .C1(KEYINPUT60), .C2(new_n826_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n303_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n826_), .ZN(G1341gat));
  AOI21_X1  g629(.A(G127gat), .B1(new_n809_), .B2(new_n614_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n585_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g632(.A(G134gat), .B1(new_n809_), .B2(new_n615_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n657_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n808_), .A2(new_n430_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n818_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n838_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT116), .B1(new_n806_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n606_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT117), .B(G141gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1344gat));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n302_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g646(.A(new_n585_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT61), .B(G155gat), .Z(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT118), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n848_), .B(new_n850_), .ZN(G1346gat));
  INV_X1    g650(.A(G162gat), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n852_), .B(new_n657_), .C1(new_n839_), .C2(new_n841_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n837_), .B1(new_n818_), .B2(new_n838_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n806_), .A2(KEYINPUT116), .A3(new_n840_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n615_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n852_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n616_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT119), .B1(new_n859_), .B2(G162gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n853_), .B1(new_n858_), .B2(new_n860_), .ZN(G1347gat));
  NOR2_X1   g660(.A1(new_n498_), .A2(new_n453_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n431_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(KEYINPUT120), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(KEYINPUT120), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n818_), .A2(new_n517_), .A3(new_n865_), .A4(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(G169gat), .B1(new_n867_), .B2(new_n606_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n866_), .ZN(new_n871_));
  NOR4_X1   g670(.A1(new_n806_), .A2(new_n377_), .A3(new_n864_), .A4(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n607_), .A3(new_n392_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n868_), .A2(new_n869_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n870_), .A2(new_n873_), .A3(new_n874_), .ZN(G1348gat));
  AOI21_X1  g674(.A(new_n389_), .B1(new_n872_), .B2(new_n302_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n867_), .A2(G176gat), .A3(new_n692_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT121), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n872_), .A2(new_n389_), .A3(new_n300_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G176gat), .B1(new_n867_), .B2(new_n303_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n882_), .ZN(G1349gat));
  OAI21_X1  g682(.A(new_n385_), .B1(new_n867_), .B2(new_n585_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n806_), .A2(new_n377_), .A3(new_n871_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n885_), .A2(new_n463_), .A3(new_n614_), .A4(new_n865_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n884_), .A2(new_n886_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1350gat));
  NAND3_X1  g689(.A1(new_n872_), .A2(new_n464_), .A3(new_n615_), .ZN(new_n891_));
  OAI21_X1  g690(.A(G190gat), .B1(new_n867_), .B2(new_n657_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1351gat));
  INV_X1    g692(.A(new_n862_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n806_), .A2(new_n430_), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n607_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n302_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n280_), .A2(KEYINPUT123), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1353gat));
  AOI21_X1  g699(.A(new_n585_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n895_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT124), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n902_), .A2(KEYINPUT126), .A3(new_n904_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n902_), .B2(new_n904_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n904_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n895_), .A2(KEYINPUT125), .A3(new_n911_), .A4(new_n901_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n907_), .A2(new_n908_), .B1(new_n910_), .B2(new_n912_), .ZN(G1354gat));
  NOR2_X1   g712(.A1(new_n806_), .A2(new_n430_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n914_), .A2(new_n615_), .A3(new_n862_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n895_), .A2(KEYINPUT127), .A3(new_n615_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n895_), .A2(G218gat), .A3(new_n658_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1355gat));
endmodule


