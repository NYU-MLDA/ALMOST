//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n963_, new_n964_, new_n966_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_, new_n980_, new_n981_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n996_,
    new_n997_, new_n998_, new_n1000_, new_n1001_, new_n1002_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1009_, new_n1010_, new_n1011_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  AOI21_X1  g005(.A(new_n205_), .B1(KEYINPUT9), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT10), .B(G99gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G106gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n207_), .A2(new_n210_), .A3(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n203_), .B(KEYINPUT6), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n218_), .A2(new_n219_), .A3(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n217_), .B1(new_n223_), .B2(new_n206_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n219_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n206_), .B1(new_n205_), .B2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(new_n216_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n215_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G64gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G57gat), .ZN(new_n230_));
  INV_X1    g029(.A(G57gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G64gat), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n230_), .A2(new_n232_), .A3(KEYINPUT11), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT67), .B(G71gat), .ZN(new_n235_));
  INV_X1    g034(.A(G78gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n235_), .A2(new_n236_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n234_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT67), .B(G71gat), .Z(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G78gat), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT11), .B1(new_n230_), .B2(new_n232_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n242_), .B(new_n237_), .C1(new_n243_), .C2(new_n233_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n228_), .A2(new_n245_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n240_), .A2(new_n244_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n223_), .A2(new_n206_), .A3(new_n217_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n226_), .A2(new_n216_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n250_), .A3(new_n215_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n246_), .A2(new_n251_), .A3(KEYINPUT12), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n228_), .A2(new_n253_), .A3(new_n245_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G230gat), .A2(G233gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n246_), .A2(new_n251_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n256_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT68), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n258_), .A2(new_n262_), .A3(new_n259_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G120gat), .B(G148gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT5), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G176gat), .B(G204gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n257_), .A2(new_n261_), .A3(new_n263_), .A4(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n262_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n271_));
  AOI211_X1 g070(.A(KEYINPUT68), .B(new_n256_), .C1(new_n246_), .C2(new_n251_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n268_), .B1(new_n273_), .B2(new_n257_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n202_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n261_), .A2(new_n263_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n259_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n267_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(KEYINPUT13), .A3(new_n269_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT69), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT37), .ZN(new_n283_));
  XOR2_X1   g082(.A(G29gat), .B(G36gat), .Z(new_n284_));
  XOR2_X1   g083(.A(G43gat), .B(G50gat), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G29gat), .B(G36gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G43gat), .B(G50gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n291_), .B(new_n215_), .C1(new_n224_), .C2(new_n227_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n210_), .A2(new_n214_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n249_), .A2(new_n248_), .B1(new_n293_), .B2(new_n207_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n290_), .B(KEYINPUT15), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n292_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT70), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT35), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n292_), .B(new_n298_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G232gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n302_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(KEYINPUT70), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT71), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G190gat), .B(G218gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(G134gat), .B(G162gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT36), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n310_), .A2(KEYINPUT36), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n306_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n313_), .ZN(new_n315_));
  AOI221_X4 g114(.A(KEYINPUT71), .B1(new_n315_), .B2(new_n311_), .C1(new_n303_), .C2(new_n305_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n283_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n306_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n303_), .A2(new_n305_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n311_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n321_), .A3(new_n315_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n316_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(KEYINPUT37), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n317_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G8gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT72), .B(G8gat), .ZN(new_n329_));
  INV_X1    g128(.A(G1gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT14), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G15gat), .B(G22gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n328_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n331_), .A2(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT73), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(new_n334_), .A3(new_n327_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G231gat), .A2(G233gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n245_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n335_), .A2(new_n336_), .A3(new_n328_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n327_), .B1(new_n339_), .B2(new_n334_), .ZN(new_n347_));
  OAI211_X1 g146(.A(G231gat), .B(G233gat), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n247_), .B1(new_n348_), .B2(new_n342_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n326_), .B1(new_n345_), .B2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G127gat), .B(G155gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT16), .ZN(new_n352_));
  XOR2_X1   g151(.A(G183gat), .B(G211gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT17), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n350_), .A2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n326_), .B(new_n356_), .C1(new_n345_), .C2(new_n349_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n354_), .ZN(new_n361_));
  OR4_X1    g160(.A1(KEYINPUT17), .A2(new_n345_), .A3(new_n349_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n325_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT75), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT99), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT18), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G64gat), .B(G92gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G169gat), .ZN(new_n372_));
  INV_X1    g171(.A(G176gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n374_), .A2(KEYINPUT24), .ZN(new_n375_));
  INV_X1    g174(.A(G183gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT25), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G183gat), .ZN(new_n379_));
  INV_X1    g178(.A(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT26), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT26), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G190gat), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n377_), .A2(new_n379_), .A3(new_n381_), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n374_), .A2(KEYINPUT24), .A3(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n375_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT76), .B(KEYINPUT23), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(new_n388_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n388_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT77), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT77), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(KEYINPUT23), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n389_), .A2(KEYINPUT76), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n396_), .B(new_n388_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n388_), .A2(KEYINPUT23), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n395_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n376_), .A2(new_n380_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT22), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G169gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n372_), .A2(KEYINPUT22), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n385_), .B1(new_n409_), .B2(G176gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n393_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G218gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G211gat), .ZN(new_n414_));
  INV_X1    g213(.A(G211gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G218gat), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT21), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G197gat), .B(G204gat), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G197gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(G204gat), .ZN(new_n422_));
  INV_X1    g221(.A(G204gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(G197gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n424_), .A3(KEYINPUT87), .ZN(new_n425_));
  OR3_X1    g224(.A1(new_n423_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n425_), .A2(KEYINPUT21), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n424_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n418_), .A2(KEYINPUT88), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT21), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n417_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT89), .B1(new_n427_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n414_), .A2(new_n416_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n419_), .B2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT21), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n420_), .B1(new_n434_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT91), .B1(new_n412_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n420_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n437_), .A2(new_n439_), .A3(new_n438_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n439_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT91), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n410_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n446_), .B(new_n447_), .C1(new_n393_), .C2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n375_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n385_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n372_), .A2(KEYINPUT79), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT78), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT22), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n453_), .A2(new_n455_), .B1(new_n407_), .B2(KEYINPUT79), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n406_), .A2(KEYINPUT78), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT79), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G169gat), .ZN(new_n459_));
  AOI21_X1  g258(.A(G176gat), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n452_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n404_), .B(new_n390_), .C1(new_n391_), .C2(new_n388_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n403_), .A2(new_n451_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n450_), .B1(new_n441_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n442_), .A2(new_n449_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G226gat), .A2(G233gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT19), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n467_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n441_), .B2(new_n463_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n403_), .A2(new_n451_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n461_), .A2(new_n462_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n446_), .A2(KEYINPUT92), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n450_), .B1(new_n412_), .B2(new_n441_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n469_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n371_), .B1(new_n468_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT27), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n465_), .A2(new_n467_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n476_), .A2(KEYINPUT93), .A3(new_n469_), .A4(new_n477_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n441_), .A2(new_n470_), .A3(new_n463_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT92), .B1(new_n446_), .B2(new_n474_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n469_), .B(new_n477_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n484_), .A2(KEYINPUT98), .A3(new_n370_), .A4(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n489_), .A2(new_n370_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT98), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n480_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n487_), .A2(new_n488_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n371_), .B1(new_n483_), .B2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT27), .B1(new_n496_), .B2(new_n491_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n498_));
  INV_X1    g297(.A(G113gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(G120gat), .ZN(new_n500_));
  INV_X1    g299(.A(G120gat), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(G113gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n498_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(G113gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(G120gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT83), .ZN(new_n506_));
  XOR2_X1   g305(.A(G127gat), .B(G134gat), .Z(new_n507_));
  NAND3_X1  g306(.A1(new_n503_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT84), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G127gat), .B(G134gat), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT83), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT83), .B1(new_n504_), .B2(new_n505_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n503_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT84), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT31), .B1(new_n510_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT84), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n512_), .A2(new_n513_), .A3(new_n511_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n507_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT31), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n509_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT82), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n388_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n401_), .B1(new_n528_), .B2(KEYINPUT77), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n387_), .B1(new_n529_), .B2(new_n400_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n457_), .A2(new_n459_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n407_), .A2(KEYINPUT79), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n458_), .B(G169gat), .C1(new_n406_), .C2(KEYINPUT78), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n373_), .A4(new_n533_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n462_), .A2(new_n534_), .A3(new_n385_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n527_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n472_), .A2(KEYINPUT30), .A3(new_n473_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(G15gat), .B(G43gat), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n536_), .A2(new_n541_), .A3(new_n537_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n526_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT82), .B1(new_n517_), .B2(new_n523_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n536_), .A2(new_n541_), .A3(new_n537_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n541_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT80), .B(KEYINPUT81), .Z(new_n548_));
  NAND2_X1  g347(.A1(G227gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G71gat), .B(G99gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n543_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G141gat), .A2(G148gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT85), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT2), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT2), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n556_), .A2(KEYINPUT85), .A3(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(G141gat), .A2(G148gat), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT3), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n558_), .A2(new_n560_), .A3(new_n563_), .A4(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G155gat), .B(G162gat), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT1), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n561_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n570_), .A2(new_n556_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n567_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n521_), .A2(new_n574_), .A3(new_n509_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n565_), .A2(new_n566_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(KEYINPUT4), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT94), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT94), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n575_), .A2(new_n577_), .A3(new_n580_), .A4(KEYINPUT4), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G225gat), .A2(G233gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n575_), .B2(KEYINPUT4), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n575_), .A2(new_n577_), .A3(new_n583_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G1gat), .B(G29gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(G85gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT0), .B(G57gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n591_), .B(new_n592_), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(new_n588_), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n585_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT97), .B1(new_n597_), .B2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n593_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n589_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n600_), .B1(new_n597_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n555_), .A2(new_n599_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n446_), .B1(new_n604_), .B2(new_n576_), .ZN(new_n605_));
  INV_X1    g404(.A(G233gat), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n606_), .A2(KEYINPUT86), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(KEYINPUT86), .ZN(new_n608_));
  OAI21_X1  g407(.A(G228gat), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n605_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G22gat), .B(G50gat), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT28), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n576_), .A2(new_n612_), .A3(new_n604_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n612_), .B1(new_n576_), .B2(new_n604_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G78gat), .B(G106gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n576_), .A2(new_n604_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT28), .ZN(new_n620_));
  INV_X1    g419(.A(new_n611_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n613_), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n616_), .A2(new_n618_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n617_), .A2(KEYINPUT90), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n616_), .B2(new_n622_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n610_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n609_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n605_), .B(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(new_n630_), .A3(new_n623_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  NOR4_X1   g431(.A1(new_n494_), .A2(new_n497_), .A3(new_n603_), .A4(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n496_), .A2(new_n491_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n575_), .A2(new_n577_), .A3(new_n584_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n600_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n575_), .A2(KEYINPUT4), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n584_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n582_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(KEYINPUT33), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n587_), .B2(new_n595_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n644_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n597_), .A2(new_n594_), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n587_), .A2(new_n589_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n596_), .A2(new_n598_), .B1(new_n649_), .B2(new_n600_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT32), .B(new_n370_), .C1(new_n468_), .C2(new_n478_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n370_), .A2(KEYINPUT32), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n489_), .A2(new_n481_), .A3(new_n482_), .A4(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  OAI22_X1  g453(.A1(new_n634_), .A2(new_n648_), .B1(new_n650_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n632_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n480_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n491_), .A2(new_n492_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n491_), .A2(new_n492_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n658_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT27), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n634_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n599_), .A2(new_n602_), .A3(new_n632_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n657_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n555_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n633_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(G229gat), .A2(G233gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n346_), .A2(new_n347_), .A3(new_n290_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n291_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n671_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n290_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n295_), .A2(new_n337_), .A3(new_n340_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n670_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(G113gat), .B(G141gat), .ZN(new_n679_));
  XNOR2_X1  g478(.A(G169gat), .B(G197gat), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n679_), .B(new_n680_), .Z(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n678_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n674_), .A2(new_n677_), .A3(new_n681_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n366_), .B1(new_n669_), .B2(new_n686_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n494_), .A2(new_n497_), .A3(new_n664_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n588_), .B1(new_n587_), .B2(new_n595_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n597_), .A2(KEYINPUT97), .A3(new_n594_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n602_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n651_), .A3(new_n653_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n587_), .A2(new_n595_), .A3(new_n644_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n646_), .B1(new_n597_), .B2(new_n594_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n496_), .A2(new_n695_), .A3(new_n491_), .A4(new_n642_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n632_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n668_), .B1(new_n688_), .B2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n494_), .A2(new_n497_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n603_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n656_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(KEYINPUT99), .A3(new_n685_), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n282_), .B(new_n365_), .C1(new_n687_), .C2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n650_), .A2(G1gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT101), .Z(new_n709_));
  NOR2_X1   g508(.A1(new_n314_), .A2(new_n316_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n280_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n685_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n363_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n702_), .A2(new_n710_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n702_), .A2(KEYINPUT102), .A3(new_n710_), .A4(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n330_), .B1(new_n719_), .B2(new_n691_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n704_), .A2(new_n707_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n705_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n709_), .A2(new_n722_), .ZN(G1324gat));
  NAND2_X1  g522(.A1(new_n661_), .A2(new_n663_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n704_), .A2(new_n329_), .A3(new_n724_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n715_), .A2(new_n699_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n727_));
  INV_X1    g526(.A(G8gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(KEYINPUT103), .B2(KEYINPUT39), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n726_), .A2(new_n727_), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n727_), .B1(new_n726_), .B2(new_n729_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n725_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT40), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(G1325gat));
  NAND2_X1  g533(.A1(new_n719_), .A2(new_n555_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G15gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT104), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n735_), .A2(new_n738_), .A3(G15gat), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT41), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G15gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n704_), .A2(new_n743_), .A3(new_n555_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n737_), .A2(KEYINPUT41), .A3(new_n739_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n744_), .A3(new_n745_), .ZN(G1326gat));
  INV_X1    g545(.A(G22gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n704_), .A2(new_n747_), .A3(new_n632_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n719_), .A2(new_n632_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G22gat), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT42), .B(new_n747_), .C1(new_n719_), .C2(new_n632_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n748_), .B(KEYINPUT105), .C1(new_n751_), .C2(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1327gat));
  NOR3_X1   g556(.A1(new_n314_), .A2(new_n283_), .A3(new_n316_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT37), .B1(new_n322_), .B2(new_n323_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n555_), .B1(new_n657_), .B2(new_n666_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n760_), .B(new_n761_), .C1(new_n762_), .C2(new_n633_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n325_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n764_));
  XOR2_X1   g563(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n712_), .A2(new_n363_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n766_), .A2(new_n767_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n650_), .ZN(new_n773_));
  INV_X1    g572(.A(G29gat), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n710_), .A2(new_n363_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n711_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n687_), .B2(new_n703_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n691_), .A2(new_n774_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT108), .ZN(new_n780_));
  OAI22_X1  g579(.A1(new_n773_), .A2(new_n774_), .B1(new_n778_), .B2(new_n780_), .ZN(G1328gat));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n782_));
  INV_X1    g581(.A(new_n776_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n699_), .A2(G36gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT99), .B1(new_n702_), .B2(new_n685_), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n366_), .B(new_n686_), .C1(new_n698_), .C2(new_n701_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n783_), .B(new_n784_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT109), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n777_), .A2(new_n789_), .A3(new_n784_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n790_), .A3(KEYINPUT45), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n771_), .A2(new_n772_), .A3(new_n699_), .ZN(new_n792_));
  INV_X1    g591(.A(G36gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT45), .B1(new_n788_), .B2(new_n790_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n782_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n795_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n772_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n766_), .A2(new_n767_), .A3(new_n770_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n724_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(G36gat), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n797_), .A2(new_n801_), .A3(KEYINPUT46), .A4(new_n791_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n796_), .A2(new_n802_), .ZN(G1329gat));
  INV_X1    g602(.A(G43gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n777_), .A2(new_n804_), .A3(new_n555_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n771_), .A2(new_n772_), .A3(new_n668_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n804_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n805_), .B(new_n808_), .C1(new_n806_), .C2(new_n804_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1330gat));
  AOI21_X1  g611(.A(G50gat), .B1(new_n777_), .B2(new_n632_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n771_), .A2(new_n772_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n632_), .A2(G50gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n813_), .B1(new_n814_), .B2(new_n815_), .ZN(G1331gat));
  NOR2_X1   g615(.A1(new_n365_), .A2(new_n711_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n669_), .A2(new_n685_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n231_), .B1(new_n819_), .B2(new_n650_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT111), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n702_), .A2(new_n710_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n363_), .A2(new_n686_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n822_), .A2(new_n281_), .A3(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n650_), .A2(new_n231_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n821_), .B1(new_n824_), .B2(new_n825_), .ZN(G1332gat));
  AOI21_X1  g625(.A(new_n229_), .B1(new_n824_), .B2(new_n724_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n819_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(new_n229_), .A3(new_n724_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1333gat));
  INV_X1    g631(.A(G71gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(new_n833_), .A3(new_n555_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n824_), .A2(new_n555_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(G71gat), .ZN(new_n837_));
  AOI211_X1 g636(.A(KEYINPUT49), .B(new_n833_), .C1(new_n824_), .C2(new_n555_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n834_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1334gat));
  NAND3_X1  g640(.A1(new_n830_), .A2(new_n236_), .A3(new_n632_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n824_), .A2(new_n632_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(G78gat), .ZN(new_n845_));
  AOI211_X1 g644(.A(KEYINPUT50), .B(new_n236_), .C1(new_n824_), .C2(new_n632_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n842_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1335gat));
  NOR3_X1   g648(.A1(new_n281_), .A2(new_n710_), .A3(new_n363_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n818_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n212_), .A3(new_n691_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n711_), .A2(new_n685_), .A3(new_n363_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n766_), .A2(new_n854_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n855_), .A2(new_n691_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n853_), .B1(new_n856_), .B2(new_n212_), .ZN(G1336gat));
  AOI21_X1  g656(.A(G92gat), .B1(new_n852_), .B2(new_n724_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n699_), .A2(new_n211_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n855_), .B2(new_n859_), .ZN(G1337gat));
  NOR3_X1   g659(.A1(new_n851_), .A2(new_n668_), .A3(new_n208_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n855_), .A2(new_n555_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(G99gat), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT51), .Z(G1338gat));
  OR3_X1    g663(.A1(new_n851_), .A2(new_n656_), .A3(new_n209_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n766_), .A2(new_n632_), .A3(new_n854_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n866_), .A2(new_n867_), .A3(G106gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n866_), .B2(G106gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n865_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g670(.A1(new_n724_), .A2(new_n632_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n668_), .A2(new_n650_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n685_), .A2(new_n269_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n252_), .A2(new_n259_), .A3(new_n254_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT55), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n877_), .A2(new_n277_), .A3(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n255_), .A2(new_n878_), .A3(new_n256_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n267_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n876_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n252_), .A2(new_n259_), .A3(new_n254_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n257_), .A2(KEYINPUT55), .A3(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n268_), .B1(new_n277_), .B2(new_n878_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n884_), .B(new_n885_), .C1(KEYINPUT116), .C2(KEYINPUT56), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n875_), .B1(new_n882_), .B2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n675_), .A2(new_n671_), .A3(new_n676_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n682_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n684_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n278_), .B2(new_n269_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n710_), .B1(new_n887_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n277_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n891_), .B1(new_n896_), .B2(new_n268_), .ZN(new_n897_));
  AND2_X1   g696(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n884_), .A2(new_n885_), .A3(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n897_), .A2(new_n899_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(KEYINPUT58), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n905_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n897_), .A2(new_n899_), .A3(new_n907_), .A4(new_n902_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n906_), .A2(new_n324_), .A3(new_n317_), .A4(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n710_), .B(KEYINPUT57), .C1(new_n887_), .C2(new_n892_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n895_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n713_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT115), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT54), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(KEYINPUT54), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n275_), .A2(new_n363_), .A3(new_n279_), .A4(new_n686_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n760_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n915_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n916_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n325_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n914_), .B1(new_n917_), .B2(new_n920_), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n912_), .A2(new_n921_), .A3(KEYINPUT119), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT119), .B1(new_n912_), .B2(new_n921_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n874_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n925_), .A2(new_n499_), .A3(new_n685_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n874_), .ZN(new_n927_));
  AOI211_X1 g726(.A(KEYINPUT59), .B(new_n927_), .C1(new_n912_), .C2(new_n921_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n928_), .B1(new_n924_), .B2(KEYINPUT59), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n929_), .A2(new_n685_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n926_), .B1(new_n930_), .B2(new_n499_), .ZN(G1340gat));
  OAI21_X1  g730(.A(new_n501_), .B1(new_n711_), .B2(KEYINPUT60), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n925_), .B(new_n932_), .C1(KEYINPUT60), .C2(new_n501_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n929_), .A2(new_n282_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n934_), .B2(new_n501_), .ZN(G1341gat));
  NAND2_X1  g734(.A1(new_n363_), .A2(G127gat), .ZN(new_n936_));
  XOR2_X1   g735(.A(new_n936_), .B(KEYINPUT120), .Z(new_n937_));
  NAND2_X1  g736(.A1(new_n929_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n925_), .A2(new_n363_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n938_), .B(KEYINPUT121), .C1(new_n940_), .C2(G127gat), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT121), .ZN(new_n942_));
  INV_X1    g741(.A(new_n937_), .ZN(new_n943_));
  AOI211_X1 g742(.A(new_n943_), .B(new_n928_), .C1(new_n924_), .C2(KEYINPUT59), .ZN(new_n944_));
  AOI21_X1  g743(.A(G127gat), .B1(new_n925_), .B2(new_n363_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n942_), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n941_), .A2(new_n946_), .ZN(G1342gat));
  INV_X1    g746(.A(G134gat), .ZN(new_n948_));
  INV_X1    g747(.A(new_n710_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n925_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n929_), .A2(new_n760_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n951_), .B2(new_n948_), .ZN(G1343gat));
  NAND2_X1  g751(.A1(new_n912_), .A2(new_n921_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n912_), .A2(new_n921_), .A3(KEYINPUT119), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n555_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n724_), .A2(new_n650_), .A3(new_n656_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n957_), .A2(new_n685_), .A3(new_n958_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g759(.A1(new_n957_), .A2(new_n282_), .A3(new_n958_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g761(.A1(new_n957_), .A2(new_n363_), .A3(new_n958_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(KEYINPUT61), .B(G155gat), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1346gat));
  NAND2_X1  g764(.A1(new_n957_), .A2(new_n958_), .ZN(new_n966_));
  OAI21_X1  g765(.A(G162gat), .B1(new_n966_), .B2(new_n325_), .ZN(new_n967_));
  OR2_X1    g766(.A1(new_n710_), .A2(G162gat), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n967_), .B1(new_n966_), .B2(new_n968_), .ZN(G1347gat));
  NAND2_X1  g768(.A1(new_n724_), .A2(new_n700_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n953_), .A2(new_n656_), .A3(new_n971_), .ZN(new_n972_));
  NOR3_X1   g771(.A1(new_n972_), .A2(new_n686_), .A3(new_n409_), .ZN(new_n973_));
  INV_X1    g772(.A(new_n972_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n372_), .B1(new_n974_), .B2(new_n685_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n973_), .B1(new_n975_), .B2(KEYINPUT62), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n976_), .B1(KEYINPUT62), .B2(new_n975_), .ZN(G1348gat));
  AOI21_X1  g776(.A(new_n632_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n978_));
  NAND4_X1  g777(.A1(new_n978_), .A2(G176gat), .A3(new_n282_), .A4(new_n971_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n373_), .B1(new_n972_), .B2(new_n711_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n980_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(KEYINPUT122), .ZN(G1349gat));
  NAND2_X1  g781(.A1(new_n377_), .A2(new_n379_), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n974_), .A2(new_n983_), .A3(new_n363_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n971_), .A2(new_n363_), .ZN(new_n985_));
  INV_X1    g784(.A(new_n985_), .ZN(new_n986_));
  OAI211_X1 g785(.A(new_n656_), .B(new_n986_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n376_), .B1(new_n987_), .B2(KEYINPUT123), .ZN(new_n988_));
  INV_X1    g787(.A(KEYINPUT123), .ZN(new_n989_));
  AOI21_X1  g788(.A(new_n989_), .B1(new_n978_), .B2(new_n986_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n984_), .B1(new_n988_), .B2(new_n990_), .ZN(new_n991_));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n991_), .A2(new_n992_), .ZN(new_n993_));
  OAI211_X1 g792(.A(KEYINPUT124), .B(new_n984_), .C1(new_n988_), .C2(new_n990_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n993_), .A2(new_n994_), .ZN(G1350gat));
  OAI21_X1  g794(.A(G190gat), .B1(new_n972_), .B2(new_n325_), .ZN(new_n996_));
  NAND3_X1  g795(.A1(new_n949_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n997_));
  XOR2_X1   g796(.A(new_n997_), .B(KEYINPUT125), .Z(new_n998_));
  OAI21_X1  g797(.A(new_n996_), .B1(new_n972_), .B2(new_n998_), .ZN(G1351gat));
  NOR2_X1   g798(.A1(new_n699_), .A2(new_n664_), .ZN(new_n1000_));
  OAI211_X1 g799(.A(new_n668_), .B(new_n1000_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n1001_));
  NOR2_X1   g800(.A1(new_n1001_), .A2(new_n686_), .ZN(new_n1002_));
  XNOR2_X1  g801(.A(new_n1002_), .B(new_n421_), .ZN(G1352gat));
  INV_X1    g802(.A(new_n1001_), .ZN(new_n1004_));
  OAI211_X1 g803(.A(new_n1004_), .B(new_n282_), .C1(KEYINPUT126), .C2(new_n423_), .ZN(new_n1005_));
  XOR2_X1   g804(.A(KEYINPUT126), .B(G204gat), .Z(new_n1006_));
  OAI21_X1  g805(.A(new_n1006_), .B1(new_n1001_), .B2(new_n281_), .ZN(new_n1007_));
  NAND2_X1  g806(.A1(new_n1005_), .A2(new_n1007_), .ZN(G1353gat));
  NOR2_X1   g807(.A1(new_n1001_), .A2(new_n713_), .ZN(new_n1009_));
  NOR3_X1   g808(.A1(new_n1009_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1010_));
  XOR2_X1   g809(.A(KEYINPUT63), .B(G211gat), .Z(new_n1011_));
  AOI21_X1  g810(.A(new_n1010_), .B1(new_n1009_), .B2(new_n1011_), .ZN(G1354gat));
  NAND3_X1  g811(.A1(new_n1004_), .A2(new_n413_), .A3(new_n949_), .ZN(new_n1013_));
  OAI21_X1  g812(.A(G218gat), .B1(new_n1001_), .B2(new_n325_), .ZN(new_n1014_));
  NAND2_X1  g813(.A1(new_n1013_), .A2(new_n1014_), .ZN(new_n1015_));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1016_));
  NAND2_X1  g815(.A1(new_n1015_), .A2(new_n1016_), .ZN(new_n1017_));
  NAND3_X1  g816(.A1(new_n1013_), .A2(new_n1014_), .A3(KEYINPUT127), .ZN(new_n1018_));
  NAND2_X1  g817(.A1(new_n1017_), .A2(new_n1018_), .ZN(G1355gat));
endmodule


