//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT77), .B(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G22gat), .ZN(new_n204_));
  INV_X1    g003(.A(G1gat), .ZN(new_n205_));
  INV_X1    g004(.A(G8gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n209_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n210_), .A2(new_n211_), .A3(new_n215_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n202_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G113gat), .B(G141gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G169gat), .B(G197gat), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n221_), .B(new_n222_), .Z(new_n223_));
  XNOR2_X1  g022(.A(new_n215_), .B(KEYINPUT15), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n212_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n212_), .A2(KEYINPUT78), .A3(new_n224_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(new_n202_), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n220_), .B(new_n223_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT79), .ZN(new_n232_));
  INV_X1    g031(.A(new_n223_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n230_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(new_n219_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n232_), .A3(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(KEYINPUT79), .B(new_n233_), .C1(new_n234_), .C2(new_n219_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240_));
  INV_X1    g039(.A(G169gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT22), .ZN(new_n242_));
  AOI21_X1  g041(.A(G176gat), .B1(new_n242_), .B2(KEYINPUT84), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(KEYINPUT84), .B2(new_n242_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT22), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G169gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT85), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n240_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT86), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G183gat), .ZN(new_n252_));
  INV_X1    g051(.A(G190gat), .ZN(new_n253_));
  OR3_X1    g052(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT23), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT23), .B1(new_n252_), .B2(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT80), .B(G190gat), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n252_), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n249_), .A2(new_n250_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G176gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n241_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n261_), .A2(new_n240_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT24), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(KEYINPUT24), .B2(new_n261_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n255_), .B(KEYINPUT83), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n264_), .B1(new_n254_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT81), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT81), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT26), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n253_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT25), .B(G183gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n257_), .A2(KEYINPUT26), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n251_), .A2(new_n259_), .B1(new_n266_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(G71gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G99gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n277_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G127gat), .B(G134gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G113gat), .B(G120gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n283_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G15gat), .B(G43gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT87), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT30), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT31), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n287_), .B(new_n291_), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G226gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT19), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n297_));
  INV_X1    g096(.A(G204gat), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n298_), .A2(G197gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(G197gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT21), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT94), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n300_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n303_), .B2(new_n299_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n301_), .B(new_n302_), .C1(new_n305_), .C2(KEYINPUT21), .ZN(new_n306_));
  INV_X1    g105(.A(new_n302_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(KEYINPUT21), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT96), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n265_), .A2(new_n254_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(G183gat), .B2(G190gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n246_), .A2(new_n242_), .A3(new_n260_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n240_), .A3(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G190gat), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n262_), .A2(new_n316_), .B1(new_n274_), .B2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n318_), .B(new_n256_), .C1(new_n261_), .C2(new_n316_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n297_), .B1(new_n311_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n309_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n277_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n296_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(new_n277_), .B2(new_n323_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n328_), .A2(KEYINPUT97), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n328_), .A2(KEYINPUT97), .B1(new_n309_), .B2(new_n320_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(new_n296_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n326_), .B1(new_n331_), .B2(KEYINPUT103), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT103), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n329_), .A2(new_n330_), .A3(new_n333_), .A4(new_n296_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G8gat), .B(G36gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G64gat), .B(G92gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT27), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n296_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n343_));
  OAI211_X1 g142(.A(KEYINPUT20), .B(new_n296_), .C1(new_n320_), .C2(new_n309_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(new_n324_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n340_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n342_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n343_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n345_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n340_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n341_), .A2(new_n348_), .B1(new_n353_), .B2(new_n342_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n323_), .B1(G228gat), .B2(G233gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(KEYINPUT1), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT89), .Z(new_n358_));
  NOR2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT88), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(KEYINPUT1), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G141gat), .A2(G148gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n360_), .A2(new_n356_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT92), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT2), .ZN(new_n372_));
  OAI22_X1  g171(.A1(new_n364_), .A2(new_n371_), .B1(new_n363_), .B2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n373_), .B1(new_n371_), .B2(new_n364_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT90), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT91), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n376_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT91), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n370_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT93), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n378_), .B(new_n379_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(KEYINPUT93), .A3(new_n370_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n367_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n355_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT95), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT95), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n390_), .B(new_n355_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G78gat), .B(G106gat), .Z(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n386_), .A2(new_n387_), .ZN(new_n395_));
  OAI211_X1 g194(.A(G228gat), .B(G233gat), .C1(new_n395_), .C2(new_n311_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n392_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n386_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT28), .B1(new_n399_), .B2(KEYINPUT29), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT28), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n386_), .A2(new_n401_), .A3(new_n387_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G22gat), .B(G50gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n400_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n406_));
  OAI22_X1  g205(.A1(new_n397_), .A2(new_n398_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n392_), .A2(new_n396_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n393_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n405_), .A2(new_n406_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n392_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT100), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n381_), .A2(new_n382_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT93), .B1(new_n384_), .B2(new_n370_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n414_), .B(new_n366_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n286_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n286_), .B1(new_n386_), .B2(new_n414_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT4), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OR3_X1    g222(.A1(new_n386_), .A2(KEYINPUT4), .A3(new_n418_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n417_), .A2(new_n418_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n386_), .A2(new_n414_), .A3(new_n286_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n422_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G85gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(KEYINPUT0), .B(G57gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n425_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n354_), .A2(new_n413_), .A3(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n425_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n351_), .A2(new_n352_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n425_), .A2(KEYINPUT33), .A3(new_n429_), .A4(new_n433_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n433_), .B1(new_n428_), .B2(new_n423_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT101), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT101), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n422_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(new_n433_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n444_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .A4(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n347_), .A2(KEYINPUT32), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n335_), .A2(new_n451_), .ZN(new_n452_));
  OR3_X1    g251(.A1(new_n343_), .A2(new_n345_), .A3(new_n451_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n452_), .B(new_n453_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n413_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n293_), .B1(new_n437_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n413_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n457_), .A2(new_n436_), .A3(new_n354_), .A4(new_n292_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n239_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT71), .ZN(new_n460_));
  INV_X1    g259(.A(G85gat), .ZN(new_n461_));
  INV_X1    g260(.A(G92gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G85gat), .A2(G92gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT9), .ZN(new_n466_));
  OR3_X1    g265(.A1(new_n465_), .A2(KEYINPUT67), .A3(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n466_), .B(new_n463_), .C1(new_n465_), .C2(KEYINPUT67), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT6), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(G99gat), .A3(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n468_), .A3(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT10), .B(G99gat), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n475_), .A2(KEYINPUT65), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(KEYINPUT65), .ZN(new_n477_));
  AOI21_X1  g276(.A(G106gat), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT66), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n479_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n474_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT8), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  INV_X1    g284(.A(G106gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n281_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n471_), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n469_), .A2(KEYINPUT6), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n484_), .B(new_n487_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n465_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n483_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n470_), .A2(new_n472_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n487_), .A2(new_n484_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT68), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT68), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n473_), .A2(new_n497_), .A3(new_n484_), .A4(new_n487_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n463_), .A2(new_n483_), .A3(new_n464_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AND4_X1   g299(.A1(KEYINPUT69), .A2(new_n496_), .A3(new_n498_), .A4(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n490_), .B2(KEYINPUT68), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT69), .B1(new_n502_), .B2(new_n498_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n493_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT70), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n496_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n502_), .A2(KEYINPUT69), .A3(new_n498_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(KEYINPUT70), .A3(new_n493_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n482_), .B1(new_n506_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G57gat), .B(G64gat), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n514_), .A2(KEYINPUT11), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G71gat), .B(G78gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(KEYINPUT11), .B2(new_n514_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n516_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT12), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n460_), .B1(new_n513_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n480_), .A2(new_n481_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n474_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT70), .B1(new_n511_), .B2(new_n493_), .ZN(new_n527_));
  AOI211_X1 g326(.A(new_n505_), .B(new_n492_), .C1(new_n509_), .C2(new_n510_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n522_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(KEYINPUT71), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n526_), .A2(new_n504_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n521_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G230gat), .A2(G233gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n536_), .B(KEYINPUT64), .Z(new_n537_));
  AOI21_X1  g336(.A(new_n482_), .B1(new_n511_), .B2(new_n493_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(new_n520_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n523_), .A2(new_n531_), .A3(new_n535_), .A4(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n520_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n533_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n537_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G120gat), .B(G148gat), .Z(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT5), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G176gat), .B(G204gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n544_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT13), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n212_), .B(new_n520_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557_));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT16), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  OR3_X1    g360(.A1(new_n556_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(KEYINPUT17), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n556_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT35), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n538_), .A2(new_n215_), .B1(new_n566_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n224_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n571_), .B1(new_n572_), .B2(new_n513_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n570_), .A2(new_n566_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI221_X1 g374(.A(new_n571_), .B1(new_n566_), .B2(new_n570_), .C1(new_n572_), .C2(new_n513_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n575_), .A2(new_n576_), .A3(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n575_), .A2(new_n576_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n579_), .B(KEYINPUT36), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT76), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n588_), .ZN(new_n589_));
  OAI221_X1 g388(.A(new_n582_), .B1(new_n587_), .B2(new_n586_), .C1(new_n583_), .C2(new_n584_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n565_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n459_), .A2(new_n553_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n436_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n205_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT38), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n585_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n553_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n599_), .A2(new_n239_), .A3(new_n565_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n205_), .B1(new_n601_), .B2(new_n593_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n596_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n595_), .B2(new_n594_), .ZN(G1324gat));
  INV_X1    g403(.A(new_n354_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n592_), .A2(new_n206_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n601_), .A2(new_n605_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n608_), .B2(G8gat), .ZN(new_n609_));
  AOI211_X1 g408(.A(KEYINPUT39), .B(new_n206_), .C1(new_n601_), .C2(new_n605_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n606_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(G1325gat));
  NAND2_X1  g412(.A1(new_n601_), .A2(new_n292_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(G15gat), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT105), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT105), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n617_), .A3(G15gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(KEYINPUT41), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(G15gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n592_), .A2(new_n620_), .A3(new_n292_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT41), .B1(new_n616_), .B2(new_n618_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1326gat));
  INV_X1    g423(.A(G22gat), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n601_), .B2(new_n413_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT42), .Z(new_n627_));
  NAND3_X1  g426(.A1(new_n592_), .A2(new_n625_), .A3(new_n413_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1327gat));
  NAND2_X1  g428(.A1(new_n597_), .A2(new_n565_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT107), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n631_), .A2(new_n553_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n459_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n593_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT44), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n589_), .A2(new_n590_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n637_), .B(KEYINPUT106), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n450_), .A2(new_n454_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n457_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n354_), .A2(new_n413_), .A3(new_n436_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n292_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n458_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n641_), .B1(new_n648_), .B2(KEYINPUT43), .ZN(new_n649_));
  INV_X1    g448(.A(new_n565_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n599_), .A2(new_n239_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n636_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n456_), .A2(new_n458_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n639_), .B1(new_n654_), .B2(new_n642_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT44), .B(new_n651_), .C1(new_n655_), .C2(new_n641_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n593_), .A2(G29gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n635_), .B1(new_n657_), .B2(new_n658_), .ZN(G1328gat));
  NAND3_X1  g458(.A1(new_n653_), .A2(new_n605_), .A3(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G36gat), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n633_), .A2(G36gat), .A3(new_n354_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT46), .B1(new_n665_), .B2(KEYINPUT108), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n667_), .B(new_n668_), .C1(new_n661_), .C2(new_n664_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n666_), .A2(new_n669_), .ZN(G1329gat));
  XNOR2_X1  g469(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n653_), .A2(new_n656_), .A3(G43gat), .A4(new_n292_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n674_));
  INV_X1    g473(.A(G43gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n675_), .B1(new_n633_), .B2(new_n293_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(new_n674_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n672_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n673_), .A2(new_n676_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT110), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n677_), .A3(new_n671_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1330gat));
  AOI21_X1  g483(.A(G50gat), .B1(new_n634_), .B2(new_n413_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n413_), .A2(G50gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n657_), .B2(new_n686_), .ZN(G1331gat));
  AOI21_X1  g486(.A(new_n238_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(new_n599_), .A3(new_n591_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G57gat), .B1(new_n689_), .B2(new_n593_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT111), .ZN(new_n691_));
  AND4_X1   g490(.A1(new_n239_), .A2(new_n598_), .A3(new_n599_), .A4(new_n650_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT112), .B(G57gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n593_), .A3(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1332gat));
  INV_X1    g494(.A(G64gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n692_), .B2(new_n605_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n689_), .A2(new_n696_), .A3(new_n605_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1333gat));
  AOI21_X1  g500(.A(new_n279_), .B1(new_n692_), .B2(new_n292_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT49), .Z(new_n703_));
  NAND2_X1  g502(.A1(new_n292_), .A2(new_n279_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT114), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n689_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1334gat));
  INV_X1    g506(.A(G78gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n692_), .B2(new_n413_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT50), .Z(new_n710_));
  NAND3_X1  g509(.A1(new_n689_), .A2(new_n708_), .A3(new_n413_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1335gat));
  AND3_X1   g511(.A1(new_n688_), .A2(new_n599_), .A3(new_n631_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n461_), .A3(new_n593_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n649_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n553_), .A2(new_n238_), .A3(new_n650_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT115), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n593_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n714_), .B1(new_n721_), .B2(new_n461_), .ZN(G1336gat));
  NAND3_X1  g521(.A1(new_n713_), .A2(new_n462_), .A3(new_n605_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n719_), .A2(new_n605_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n723_), .B1(new_n725_), .B2(new_n462_), .ZN(G1337gat));
  OAI21_X1  g525(.A(G99gat), .B1(new_n718_), .B2(new_n293_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n476_), .A2(new_n477_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n713_), .A2(new_n292_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g530(.A1(new_n713_), .A2(new_n486_), .A3(new_n413_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n413_), .B(new_n717_), .C1(new_n655_), .C2(new_n641_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(G106gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n733_), .B2(G106gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g537(.A1(new_n217_), .A2(new_n218_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n223_), .B1(new_n739_), .B2(new_n202_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n218_), .A2(G229gat), .A3(G233gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(new_n229_), .B2(new_n741_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n231_), .A2(KEYINPUT117), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT117), .B1(new_n231_), .B2(new_n742_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n544_), .A2(new_n548_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n523_), .A2(new_n531_), .A3(new_n535_), .A4(new_n541_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n537_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n540_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n534_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n532_), .B2(new_n521_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n529_), .A2(new_n530_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n460_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n755_), .A2(KEYINPUT55), .A3(new_n531_), .A4(new_n539_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n749_), .A2(new_n751_), .A3(new_n756_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n548_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT56), .B1(new_n757_), .B2(new_n548_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n747_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n747_), .B(KEYINPUT58), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n638_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n746_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n238_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n757_), .A2(new_n548_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n548_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n551_), .A2(new_n745_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT57), .B(new_n585_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n764_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n585_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(new_n650_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n553_), .A2(new_n591_), .A3(new_n239_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n778_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n457_), .A2(new_n354_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n593_), .A2(new_n292_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OR3_X1    g585(.A1(new_n782_), .A2(KEYINPUT59), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n765_), .A2(new_n238_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n772_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n597_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n792_), .B2(KEYINPUT57), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n776_), .A2(KEYINPUT118), .A3(new_n775_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n773_), .A4(new_n764_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n781_), .B1(new_n795_), .B2(new_n565_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT59), .B1(new_n796_), .B2(new_n786_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n787_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(G113gat), .B1(new_n798_), .B2(new_n239_), .ZN(new_n799_));
  OR3_X1    g598(.A1(new_n796_), .A2(KEYINPUT119), .A3(new_n786_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT119), .B1(new_n796_), .B2(new_n786_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(G113gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n238_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n799_), .A2(new_n804_), .ZN(G1340gat));
  OAI21_X1  g604(.A(G120gat), .B1(new_n798_), .B2(new_n553_), .ZN(new_n806_));
  INV_X1    g605(.A(G120gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n553_), .B2(KEYINPUT60), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n802_), .B(new_n808_), .C1(KEYINPUT60), .C2(new_n807_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n809_), .ZN(G1341gat));
  OAI21_X1  g609(.A(G127gat), .B1(new_n798_), .B2(new_n565_), .ZN(new_n811_));
  INV_X1    g610(.A(G127gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n802_), .A2(new_n812_), .A3(new_n650_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1342gat));
  NAND3_X1  g613(.A1(new_n800_), .A2(new_n597_), .A3(new_n801_), .ZN(new_n815_));
  INV_X1    g614(.A(G134gat), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(KEYINPUT120), .A3(new_n816_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n787_), .A2(new_n797_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(KEYINPUT121), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n816_), .A2(KEYINPUT121), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n637_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n819_), .A2(new_n820_), .B1(new_n821_), .B2(new_n824_), .ZN(G1343gat));
  NOR4_X1   g624(.A1(new_n605_), .A2(new_n457_), .A3(new_n436_), .A4(new_n292_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT118), .B1(new_n776_), .B2(new_n775_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n774_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n650_), .B1(new_n828_), .B2(new_n794_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT122), .B(new_n826_), .C1(new_n829_), .C2(new_n781_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  INV_X1    g630(.A(new_n826_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n796_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n238_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n599_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n650_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT61), .B(G155gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1346gat));
  INV_X1    g640(.A(G162gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n834_), .B2(new_n642_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n585_), .A2(G162gat), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT123), .B1(new_n843_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n846_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n849_));
  INV_X1    g648(.A(new_n642_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n848_), .B(new_n849_), .C1(new_n842_), .C2(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n847_), .A2(new_n852_), .ZN(G1347gat));
  NAND2_X1  g652(.A1(new_n436_), .A2(new_n292_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n354_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n457_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n782_), .A2(new_n239_), .A3(new_n856_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n858_));
  OR3_X1    g657(.A1(new_n857_), .A2(new_n241_), .A3(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n857_), .B2(new_n241_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n857_), .A2(new_n246_), .A3(new_n242_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(G1348gat));
  NOR2_X1   g661(.A1(new_n782_), .A2(new_n856_), .ZN(new_n863_));
  AOI21_X1  g662(.A(G176gat), .B1(new_n863_), .B2(new_n599_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n796_), .A2(new_n413_), .ZN(new_n865_));
  NOR4_X1   g664(.A1(new_n553_), .A2(new_n854_), .A3(new_n260_), .A4(new_n354_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(G1349gat));
  INV_X1    g666(.A(new_n863_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n868_), .A2(new_n274_), .A3(new_n565_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n865_), .A2(new_n650_), .A3(new_n855_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(G183gat), .B1(new_n870_), .B2(new_n871_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n869_), .B1(new_n872_), .B2(new_n873_), .ZN(G1350gat));
  OAI21_X1  g673(.A(G190gat), .B1(new_n868_), .B2(new_n637_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n863_), .A2(new_n317_), .A3(new_n597_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1351gat));
  NAND3_X1  g676(.A1(new_n413_), .A2(new_n436_), .A3(new_n293_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n796_), .A2(new_n354_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n238_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g680(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT126), .B(G204gat), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n599_), .ZN(new_n884_));
  MUX2_X1   g683(.A(new_n882_), .B(new_n883_), .S(new_n884_), .Z(G1353gat));
  NAND2_X1  g684(.A1(new_n879_), .A2(new_n650_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n887_));
  AND2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(new_n886_), .B2(new_n887_), .ZN(G1354gat));
  NAND2_X1  g689(.A1(new_n879_), .A2(new_n597_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT127), .B(G218gat), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n637_), .A2(new_n892_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n891_), .A2(new_n892_), .B1(new_n879_), .B2(new_n893_), .ZN(G1355gat));
endmodule


