//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n203_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n210_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT80), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(G169gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n204_), .A2(KEYINPUT22), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n205_), .A3(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n216_), .B1(new_n217_), .B2(G169gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n208_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT81), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n222_), .A2(new_n223_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n215_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G227gat), .A2(G233gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n229_), .B(KEYINPUT82), .Z(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n228_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G71gat), .B(G99gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n235_), .A2(KEYINPUT83), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(KEYINPUT83), .ZN(new_n237_));
  XOR2_X1   g036(.A(G113gat), .B(G120gat), .Z(new_n238_));
  OR3_X1    g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n238_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT31), .ZN(new_n242_));
  XOR2_X1   g041(.A(G15gat), .B(G43gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n234_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n234_), .A2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(G155gat), .A2(G162gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249_));
  INV_X1    g048(.A(G141gat), .ZN(new_n250_));
  INV_X1    g049(.A(G148gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT84), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n252_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT2), .Z(new_n257_));
  OAI211_X1 g056(.A(new_n248_), .B(new_n249_), .C1(new_n255_), .C2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n249_), .A2(KEYINPUT1), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n248_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n249_), .A2(KEYINPUT1), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n252_), .B(new_n256_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n241_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n239_), .A2(new_n258_), .A3(new_n262_), .A4(new_n240_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G225gat), .A2(G233gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(KEYINPUT4), .A3(new_n265_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n241_), .A2(new_n271_), .A3(new_n263_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n267_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G1gat), .B(G29gat), .ZN(new_n274_));
  INV_X1    g073(.A(G85gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT0), .B(G57gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n269_), .A2(new_n273_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT98), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n269_), .B2(new_n273_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(KEYINPUT98), .B(new_n278_), .C1(new_n269_), .C2(new_n273_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n247_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n263_), .A2(KEYINPUT29), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT86), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n286_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G22gat), .B(G50gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G228gat), .A2(G233gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n263_), .A2(KEYINPUT29), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT88), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT89), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G204gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT90), .B1(new_n297_), .B2(G197gat), .ZN(new_n298_));
  INV_X1    g097(.A(G197gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(G204gat), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n297_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT21), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT91), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n297_), .B2(G197gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n299_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n305_), .B(new_n306_), .C1(new_n299_), .C2(G204gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n302_), .B(new_n303_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n303_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(KEYINPUT21), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n293_), .B1(new_n296_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT89), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT88), .B1(new_n293_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n294_), .A2(new_n312_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G78gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n314_), .A2(G78gat), .A3(new_n317_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(G106gat), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT87), .ZN(new_n323_));
  AOI21_X1  g122(.A(G106gat), .B1(new_n320_), .B2(new_n321_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n292_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n321_), .ZN(new_n326_));
  INV_X1    g125(.A(G106gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n328_), .A2(KEYINPUT87), .A3(new_n291_), .A4(new_n322_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT19), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT93), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n211_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n213_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n208_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT22), .B(G169gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n205_), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n335_), .A2(new_n210_), .B1(new_n225_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT20), .B1(new_n313_), .B2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n228_), .A2(new_n312_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n332_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G8gat), .B(G36gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT18), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n228_), .A2(new_n312_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n313_), .A2(new_n339_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n332_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT20), .A4(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n342_), .A2(new_n346_), .A3(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n340_), .A2(new_n341_), .A3(new_n332_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n211_), .B(KEYINPUT93), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n210_), .B1(new_n353_), .B2(new_n214_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n225_), .A2(new_n338_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT20), .B1(new_n356_), .B2(new_n312_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n357_), .A2(KEYINPUT97), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(KEYINPUT97), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n347_), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n352_), .B1(new_n360_), .B2(new_n332_), .ZN(new_n361_));
  OAI211_X1 g160(.A(KEYINPUT27), .B(new_n351_), .C1(new_n361_), .C2(new_n346_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n346_), .B1(new_n342_), .B2(new_n350_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT94), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(new_n351_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n351_), .A2(new_n364_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT27), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT100), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI211_X1 g168(.A(KEYINPUT100), .B(KEYINPUT27), .C1(new_n365_), .C2(new_n366_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n330_), .B(new_n362_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT102), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n367_), .B(new_n368_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n374_), .A2(KEYINPUT102), .A3(new_n330_), .A4(new_n362_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n285_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n247_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n281_), .A2(KEYINPUT33), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT33), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n379_), .B(new_n278_), .C1(new_n269_), .C2(new_n273_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n278_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n270_), .A2(KEYINPUT95), .A3(new_n267_), .A4(new_n272_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n270_), .A2(new_n267_), .A3(new_n272_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT95), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n365_), .A2(new_n366_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT96), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n378_), .A2(new_n380_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT96), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n366_), .A4(new_n365_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n361_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n342_), .A2(new_n350_), .A3(new_n395_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n396_), .A2(new_n282_), .A3(new_n283_), .A4(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n391_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n330_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT99), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n325_), .A2(new_n284_), .A3(new_n329_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n402_), .A2(new_n374_), .A3(KEYINPUT101), .A4(new_n362_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT101), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n362_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n325_), .A2(new_n284_), .A3(new_n329_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT99), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n399_), .A2(new_n408_), .A3(new_n330_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n401_), .A2(new_n403_), .A3(new_n407_), .A4(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n376_), .B1(new_n377_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G29gat), .B(G36gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G43gat), .B(G50gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT76), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G15gat), .B(G22gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G1gat), .A2(G8gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT14), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G1gat), .B(G8gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n415_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT77), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n415_), .A2(new_n422_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT78), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G229gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n414_), .B(KEYINPUT15), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n422_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n425_), .A2(new_n430_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G113gat), .B(G141gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G169gat), .B(G197gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  NOR2_X1   g238(.A1(new_n439_), .A2(KEYINPUT79), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n440_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n411_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G231gat), .A2(G233gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n421_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G57gat), .B(G64gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G71gat), .B(G78gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT11), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  INV_X1    g249(.A(G64gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G57gat), .ZN(new_n452_));
  INV_X1    g251(.A(G57gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G64gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n454_), .A3(KEYINPUT11), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n447_), .A2(KEYINPUT11), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n449_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n446_), .B(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G127gat), .B(G155gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT16), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G183gat), .B(G211gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT17), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n459_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT75), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n463_), .A2(new_n464_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n459_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G230gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(G92gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n275_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT6), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT7), .ZN(new_n483_));
  INV_X1    g282(.A(G99gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n327_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n477_), .B1(new_n482_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT8), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n480_), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n478_), .A2(KEYINPUT6), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n486_), .B(new_n485_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n477_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT64), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n496_), .A2(KEYINPUT9), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(KEYINPUT9), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n497_), .A2(G85gat), .A3(G92gat), .A4(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n474_), .A2(new_n496_), .A3(KEYINPUT9), .A4(new_n475_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n479_), .A2(new_n481_), .ZN(new_n501_));
  OR2_X1    g300(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n327_), .A3(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .A4(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n458_), .B1(new_n495_), .B2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(KEYINPUT65), .ZN(new_n507_));
  INV_X1    g306(.A(new_n486_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  AOI211_X1 g309(.A(KEYINPUT8), .B(new_n476_), .C1(new_n510_), .C2(new_n501_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n493_), .B1(new_n492_), .B2(new_n477_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n505_), .B(new_n458_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n472_), .B1(new_n507_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(new_n513_), .B2(new_n507_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n513_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n516_), .B1(KEYINPUT12), .B2(new_n506_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT66), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n505_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n458_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT12), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n518_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AOI211_X1 g322(.A(KEYINPUT66), .B(KEYINPUT12), .C1(new_n519_), .C2(new_n520_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n517_), .B(new_n472_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n515_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G120gat), .B(G148gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(G176gat), .B(G204gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n526_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n526_), .A2(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT13), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n537_), .B(KEYINPUT68), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n540_));
  NOR2_X1   g339(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n541_));
  INV_X1    g340(.A(new_n505_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n414_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT71), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n543_), .A2(KEYINPUT71), .A3(new_n414_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n433_), .A2(new_n519_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OR3_X1    g354(.A1(new_n549_), .A2(KEYINPUT72), .A3(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT73), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n549_), .A2(new_n550_), .B1(KEYINPUT36), .B2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n555_), .B1(new_n549_), .B2(KEYINPUT72), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n560_), .A2(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n556_), .A2(new_n561_), .A3(new_n566_), .A4(new_n562_), .ZN(new_n567_));
  AOI211_X1 g366(.A(new_n540_), .B(new_n541_), .C1(new_n565_), .C2(new_n567_), .ZN(new_n568_));
  AND4_X1   g367(.A1(KEYINPUT74), .A2(new_n565_), .A3(KEYINPUT37), .A4(new_n567_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n444_), .A2(new_n471_), .A3(new_n539_), .A4(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n571_), .A2(G1gat), .A3(new_n284_), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n572_), .B(KEYINPUT38), .Z(new_n573_));
  INV_X1    g372(.A(KEYINPUT104), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n410_), .A2(new_n377_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n376_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n565_), .A2(new_n567_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n574_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n411_), .A2(KEYINPUT104), .A3(new_n578_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n441_), .A2(new_n442_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n537_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT103), .Z(new_n585_));
  AND2_X1   g384(.A1(new_n585_), .A2(new_n471_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n284_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(G1gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n573_), .A2(new_n590_), .ZN(G1324gat));
  OAI211_X1 g390(.A(new_n405_), .B(new_n586_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(KEYINPUT106), .A3(G8gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT39), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT106), .B1(new_n592_), .B2(G8gat), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n405_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(G8gat), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OR3_X1    g400(.A1(new_n571_), .A2(KEYINPUT105), .A3(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT105), .B1(new_n571_), .B2(new_n601_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OR3_X1    g406(.A1(new_n596_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n607_), .B1(new_n596_), .B2(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(G1325gat));
  INV_X1    g409(.A(G15gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n587_), .B2(new_n247_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(KEYINPUT41), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(KEYINPUT41), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n247_), .A2(new_n611_), .ZN(new_n615_));
  OAI22_X1  g414(.A1(new_n613_), .A2(new_n614_), .B1(new_n571_), .B2(new_n615_), .ZN(G1326gat));
  INV_X1    g415(.A(G22gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n330_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n587_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT42), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(new_n620_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n618_), .A2(new_n617_), .ZN(new_n623_));
  OAI22_X1  g422(.A1(new_n621_), .A2(new_n622_), .B1(new_n571_), .B2(new_n623_), .ZN(G1327gat));
  NOR2_X1   g423(.A1(new_n471_), .A2(new_n579_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(new_n537_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n444_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G29gat), .B1(new_n628_), .B2(new_n588_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n585_), .A2(new_n470_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT43), .B1(new_n570_), .B2(KEYINPUT108), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(new_n411_), .B2(new_n570_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n570_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n403_), .A2(new_n407_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n399_), .A2(new_n408_), .A3(new_n330_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n408_), .B1(new_n399_), .B2(new_n330_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n247_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n634_), .B(new_n631_), .C1(new_n639_), .C2(new_n376_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n630_), .B1(new_n633_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT44), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n642_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n588_), .A2(G29gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n629_), .B1(new_n645_), .B2(new_n646_), .ZN(G1328gat));
  NOR2_X1   g446(.A1(new_n599_), .A2(G36gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n627_), .A2(KEYINPUT110), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT110), .B1(new_n627_), .B2(new_n649_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(KEYINPUT45), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT45), .B1(new_n650_), .B2(new_n651_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G36gat), .B1(new_n644_), .B2(new_n599_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n654_), .A2(KEYINPUT46), .A3(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1329gat));
  NAND3_X1  g459(.A1(new_n645_), .A2(G43gat), .A3(new_n247_), .ZN(new_n661_));
  INV_X1    g460(.A(G43gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n627_), .B2(new_n377_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT47), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(new_n666_), .A3(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1330gat));
  OR3_X1    g467(.A1(new_n627_), .A2(G50gat), .A3(new_n330_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n645_), .A2(KEYINPUT111), .A3(new_n618_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G50gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT111), .B1(new_n645_), .B2(new_n618_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n669_), .B1(new_n671_), .B2(new_n672_), .ZN(G1331gat));
  NOR2_X1   g472(.A1(new_n411_), .A2(new_n583_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n634_), .A2(new_n470_), .A3(new_n537_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n453_), .B1(new_n676_), .B2(new_n284_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT112), .Z(new_n678_));
  NOR2_X1   g477(.A1(new_n583_), .A2(new_n470_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n582_), .A2(new_n538_), .A3(new_n679_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n680_), .A2(new_n453_), .A3(new_n284_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n678_), .A2(new_n681_), .ZN(G1332gat));
  INV_X1    g481(.A(new_n676_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n451_), .A3(new_n405_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G64gat), .B1(new_n680_), .B2(new_n599_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(KEYINPUT48), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(KEYINPUT48), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(new_n686_), .B2(new_n687_), .ZN(G1333gat));
  OR3_X1    g487(.A1(new_n676_), .A2(G71gat), .A3(new_n377_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G71gat), .B1(new_n680_), .B2(new_n377_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(KEYINPUT49), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(KEYINPUT49), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(G1334gat));
  NAND3_X1  g492(.A1(new_n683_), .A2(new_n319_), .A3(new_n618_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G78gat), .B1(new_n680_), .B2(new_n330_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT50), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT50), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(G1335gat));
  NOR3_X1   g497(.A1(new_n537_), .A2(new_n471_), .A3(new_n583_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n633_), .B2(new_n640_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G85gat), .B1(new_n702_), .B2(new_n284_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n674_), .A2(new_n538_), .A3(new_n625_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n588_), .A2(new_n275_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(G1336gat));
  OAI21_X1  g505(.A(G92gat), .B1(new_n702_), .B2(new_n599_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n405_), .A2(new_n473_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n704_), .B2(new_n708_), .ZN(G1337gat));
  OAI21_X1  g508(.A(G99gat), .B1(new_n702_), .B2(new_n377_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n247_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n704_), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g512(.A(new_n327_), .B1(new_n701_), .B2(new_n618_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT52), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT115), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n631_), .B1(new_n577_), .B2(new_n634_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n411_), .A2(new_n570_), .A3(new_n632_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n618_), .B(new_n699_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n715_), .A3(G106gat), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT114), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(G106gat), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT115), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(KEYINPUT52), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n714_), .A2(KEYINPUT114), .A3(new_n715_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n716_), .A2(new_n722_), .A3(new_n725_), .A4(new_n726_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n704_), .A2(G106gat), .A3(new_n330_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT113), .Z(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT53), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT53), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n727_), .A2(new_n732_), .A3(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1339gat));
  NAND2_X1  g533(.A1(new_n373_), .A2(new_n375_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n377_), .A2(new_n284_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n432_), .A2(new_n439_), .A3(new_n435_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n429_), .A2(new_n431_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n430_), .B1(new_n425_), .B2(new_n434_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n738_), .B1(new_n741_), .B2(new_n439_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(new_n533_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n517_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n472_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(KEYINPUT55), .A3(new_n525_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n519_), .A2(KEYINPUT12), .A3(new_n520_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n513_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT66), .B1(new_n506_), .B2(KEYINPUT12), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n521_), .A2(new_n518_), .A3(new_n522_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n472_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n747_), .A2(KEYINPUT117), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT117), .B1(new_n747_), .B2(new_n754_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  NOR4_X1   g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .A4(new_n531_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n747_), .A2(new_n754_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n531_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n747_), .A2(KEYINPUT117), .A3(new_n754_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT56), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n743_), .B1(new_n758_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT58), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n570_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n759_), .A2(new_n760_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n532_), .A3(new_n762_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n757_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n761_), .A2(KEYINPUT56), .A3(new_n762_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n771_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n743_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT58), .B(new_n743_), .C1(new_n758_), .C2(new_n763_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n766_), .A2(new_n772_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n583_), .A2(new_n534_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n770_), .B1(new_n763_), .B2(KEYINPUT118), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n755_), .A2(new_n756_), .A3(new_n531_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(KEYINPUT56), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n742_), .B1(new_n535_), .B2(new_n534_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n578_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n776_), .B1(new_n786_), .B2(KEYINPUT57), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n781_), .B1(new_n780_), .B2(KEYINPUT56), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n768_), .A2(KEYINPUT118), .A3(new_n757_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n770_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n784_), .B1(new_n790_), .B2(new_n778_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n578_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n470_), .B1(new_n787_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n537_), .A2(new_n679_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT116), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n537_), .A2(new_n679_), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n634_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n737_), .B1(new_n794_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(G113gat), .B1(new_n802_), .B2(new_n583_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n737_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(KEYINPUT120), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n737_), .B2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n805_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT121), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n794_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n792_), .B1(new_n791_), .B2(new_n578_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n758_), .B1(new_n781_), .B2(new_n769_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n777_), .B1(new_n814_), .B2(new_n789_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n579_), .C1(new_n815_), .C2(new_n784_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n816_), .A3(new_n776_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(KEYINPUT121), .A3(new_n470_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n812_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n810_), .B1(new_n819_), .B2(new_n801_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n794_), .A2(new_n801_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n804_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n820_), .B1(KEYINPUT59), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n583_), .A2(G113gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT122), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n803_), .B1(new_n823_), .B2(new_n825_), .ZN(G1340gat));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n538_), .B1(new_n802_), .B2(new_n806_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n820_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n539_), .B1(new_n822_), .B2(KEYINPUT59), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n817_), .A2(KEYINPUT121), .A3(new_n470_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT121), .B1(new_n817_), .B2(new_n470_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n801_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n809_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(new_n834_), .A3(KEYINPUT123), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n829_), .A2(new_n835_), .A3(G120gat), .ZN(new_n836_));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n537_), .B2(KEYINPUT60), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n802_), .B(new_n838_), .C1(KEYINPUT60), .C2(new_n837_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT124), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT124), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n836_), .A2(new_n842_), .A3(new_n839_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n802_), .B2(new_n471_), .ZN(new_n845_));
  INV_X1    g644(.A(G127gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n471_), .B2(KEYINPUT125), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(KEYINPUT125), .B2(new_n846_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n845_), .B1(new_n823_), .B2(new_n848_), .ZN(G1342gat));
  INV_X1    g648(.A(G134gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n802_), .A2(new_n850_), .A3(new_n578_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n823_), .A2(new_n634_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n853_), .B2(new_n850_), .ZN(G1343gat));
  NOR4_X1   g653(.A1(new_n405_), .A2(new_n330_), .A3(new_n284_), .A4(new_n247_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n821_), .A2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT126), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n443_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n250_), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n539_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n251_), .ZN(G1345gat));
  NOR2_X1   g660(.A1(new_n857_), .A2(new_n470_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT61), .B(G155gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  OAI21_X1  g663(.A(G162gat), .B1(new_n857_), .B2(new_n570_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n579_), .A2(G162gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n857_), .B2(new_n866_), .ZN(G1347gat));
  AOI21_X1  g666(.A(new_n204_), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n599_), .A2(new_n285_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n618_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n833_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n872_), .B2(new_n443_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n443_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n873_), .A2(new_n874_), .B1(new_n875_), .B2(new_n337_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n873_), .B2(new_n874_), .ZN(G1348gat));
  OR2_X1    g676(.A1(new_n872_), .A2(new_n537_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n821_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n618_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n539_), .A2(new_n205_), .A3(new_n870_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n878_), .A2(new_n205_), .B1(new_n880_), .B2(new_n881_), .ZN(G1349gat));
  NOR2_X1   g681(.A1(new_n870_), .A2(new_n470_), .ZN(new_n883_));
  AOI21_X1  g682(.A(G183gat), .B1(new_n880_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n872_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n471_), .A2(new_n353_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n884_), .B1(new_n885_), .B2(new_n887_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n872_), .B2(new_n570_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n578_), .A2(new_n213_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n872_), .B2(new_n890_), .ZN(G1351gat));
  NOR4_X1   g690(.A1(new_n879_), .A2(new_n247_), .A3(new_n599_), .A4(new_n406_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n583_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n538_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g695(.A1(new_n892_), .A2(new_n471_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  AND2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n897_), .B2(new_n898_), .ZN(G1354gat));
  INV_X1    g700(.A(G218gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n892_), .A2(new_n902_), .A3(new_n578_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n892_), .A2(new_n634_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n902_), .ZN(G1355gat));
endmodule


