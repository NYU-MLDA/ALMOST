//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND4_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(G183gat), .A4(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT23), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n203_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n204_), .B1(new_n208_), .B2(new_n202_), .ZN(new_n209_));
  NOR3_X1   g008(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT25), .B(G183gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n214_), .A2(new_n218_), .A3(KEYINPUT91), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT91), .B1(new_n214_), .B2(new_n218_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n211_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G218gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n222_), .A2(G211gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(G211gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT87), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G211gat), .B(G218gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT87), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G197gat), .B(G204gat), .Z(new_n229_));
  NAND4_X1  g028(.A1(new_n225_), .A2(new_n228_), .A3(KEYINPUT21), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(KEYINPUT21), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G197gat), .B(G204gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT21), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n226_), .A2(new_n227_), .ZN(new_n235_));
  NOR3_X1   g034(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT87), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n231_), .B(new_n234_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G169gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n208_), .ZN(new_n240_));
  OR2_X1    g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n239_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n221_), .A2(new_n230_), .A3(new_n237_), .A4(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n239_), .B1(new_n209_), .B2(new_n242_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n246_));
  INV_X1    g045(.A(G190gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT26), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n247_), .A2(KEYINPUT26), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n212_), .B(new_n248_), .C1(new_n249_), .C2(new_n246_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n210_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n216_), .A2(KEYINPUT82), .A3(new_n217_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT82), .B1(new_n216_), .B2(new_n217_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n250_), .B(new_n251_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n245_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n237_), .A2(new_n230_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n244_), .A2(KEYINPUT20), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G226gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT19), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT96), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT20), .B1(new_n255_), .B2(new_n256_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT90), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n221_), .A2(new_n243_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n264_), .A2(new_n265_), .B1(new_n266_), .B2(new_n256_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n260_), .ZN(new_n268_));
  OAI211_X1 g067(.A(KEYINPUT90), .B(KEYINPUT20), .C1(new_n255_), .C2(new_n256_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n258_), .A2(KEYINPUT96), .A3(new_n260_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n263_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G8gat), .B(G36gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT18), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT99), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  AND4_X1   g077(.A1(KEYINPUT20), .A2(new_n244_), .A3(new_n268_), .A4(new_n257_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n264_), .A2(new_n265_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n266_), .A2(new_n256_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n269_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n260_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n276_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n278_), .A2(KEYINPUT27), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n268_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n276_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n287_), .A2(new_n279_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(new_n260_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n279_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n276_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n286_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n285_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT2), .ZN(new_n296_));
  INV_X1    g095(.A(G141gat), .ZN(new_n297_));
  INV_X1    g096(.A(G148gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n299_), .A2(new_n301_), .A3(new_n302_), .A4(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(KEYINPUT1), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(G155gat), .A3(G162gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n311_), .A3(new_n305_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G141gat), .B(G148gat), .Z(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT29), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n256_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G228gat), .ZN(new_n318_));
  INV_X1    g117(.A(G233gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n320_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n256_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G78gat), .B(G106gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(KEYINPUT88), .ZN(new_n328_));
  INV_X1    g127(.A(new_n323_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n322_), .B1(new_n256_), .B2(new_n316_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n324_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT88), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(new_n315_), .B2(KEYINPUT29), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n304_), .A2(new_n307_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337_));
  INV_X1    g136(.A(new_n334_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G22gat), .B(G50gat), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n335_), .A2(new_n341_), .A3(new_n339_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT86), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT86), .B1(new_n343_), .B2(new_n344_), .ZN(new_n348_));
  OAI22_X1  g147(.A1(new_n328_), .A2(new_n333_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n331_), .A2(new_n345_), .A3(new_n326_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n349_), .A2(KEYINPUT89), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT89), .B1(new_n349_), .B2(new_n350_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n295_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G227gat), .A2(G233gat), .ZN(new_n355_));
  INV_X1    g154(.A(G71gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G99gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n255_), .B(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G127gat), .B(G134gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(G113gat), .B(G120gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  XNOR2_X1  g161(.A(new_n359_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G15gat), .B(G43gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT84), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT30), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT31), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n363_), .B(new_n367_), .Z(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n336_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n362_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n360_), .B(new_n361_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n372_), .A3(new_n336_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n371_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n362_), .A2(KEYINPUT4), .A3(new_n336_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n370_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n369_), .A3(new_n376_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT97), .B1(new_n381_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT97), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n379_), .A2(new_n380_), .A3(new_n389_), .A4(new_n386_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n368_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n354_), .A2(new_n395_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n379_), .A2(new_n380_), .A3(new_n386_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n391_), .B1(new_n397_), .B2(new_n389_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n276_), .A2(KEYINPUT32), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n398_), .A2(new_n388_), .B1(new_n272_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n290_), .A2(new_n291_), .A3(new_n399_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT95), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT95), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n283_), .A2(new_n404_), .A3(new_n399_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n374_), .A2(new_n376_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n378_), .B1(new_n407_), .B2(KEYINPUT4), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT94), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n369_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n387_), .B1(new_n370_), .B2(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n409_), .B1(new_n408_), .B2(new_n369_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT33), .B1(new_n381_), .B2(new_n387_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT33), .ZN(new_n416_));
  AOI211_X1 g215(.A(new_n416_), .B(new_n386_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n289_), .A2(new_n292_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n401_), .A2(new_n406_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n352_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n349_), .A2(KEYINPUT89), .A3(new_n350_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT98), .B1(new_n420_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n272_), .A2(new_n400_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n404_), .B1(new_n283_), .B2(new_n399_), .ZN(new_n426_));
  NOR4_X1   g225(.A1(new_n287_), .A2(KEYINPUT95), .A3(new_n279_), .A4(new_n400_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n393_), .B(new_n425_), .C1(new_n426_), .C2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n415_), .A2(new_n417_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n412_), .A2(new_n413_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n288_), .B1(new_n287_), .B2(new_n279_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n284_), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT98), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n353_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n295_), .A2(new_n423_), .A3(new_n394_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n424_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n368_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n396_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(G230gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n319_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT64), .ZN(new_n444_));
  NAND2_X1  g243(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n445_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT64), .B1(new_n447_), .B2(new_n442_), .ZN(new_n448_));
  AOI21_X1  g247(.A(G106gat), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G99gat), .A2(G106gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT6), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(G99gat), .A3(G106gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G85gat), .ZN(new_n455_));
  INV_X1    g254(.A(G92gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G85gat), .A2(G92gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(KEYINPUT9), .A3(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n454_), .B(new_n459_), .C1(KEYINPUT9), .C2(new_n458_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n449_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT65), .ZN(new_n462_));
  OAI221_X1 g261(.A(new_n462_), .B1(KEYINPUT66), .B2(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G99gat), .A2(G106gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n465_), .B2(KEYINPUT65), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT7), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT65), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n454_), .A2(new_n463_), .A3(new_n466_), .A4(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n457_), .A2(new_n458_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT8), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n473_), .A2(KEYINPUT68), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT67), .B1(new_n473_), .B2(KEYINPUT68), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n477_), .B1(KEYINPUT67), .B2(new_n473_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n469_), .A2(new_n471_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n461_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G57gat), .B(G64gat), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n483_));
  XOR2_X1   g282(.A(G71gat), .B(G78gat), .Z(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n483_), .A2(new_n484_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n480_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n480_), .A2(new_n487_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n441_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(new_n480_), .B2(new_n487_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT69), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n469_), .A2(new_n471_), .A3(new_n478_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n474_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n463_), .A2(new_n466_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n451_), .A2(new_n453_), .B1(KEYINPUT65), .B2(new_n467_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n470_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT69), .B(new_n479_), .C1(new_n500_), .C2(new_n474_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n461_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n485_), .A2(KEYINPUT12), .A3(new_n486_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n493_), .B(new_n488_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n491_), .B1(new_n504_), .B2(new_n441_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G120gat), .B(G148gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT5), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G176gat), .B(G204gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n509_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT13), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(KEYINPUT13), .A3(new_n511_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G29gat), .B(G36gat), .Z(new_n518_));
  XOR2_X1   g317(.A(G43gat), .B(G50gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT15), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT75), .B(G8gat), .ZN(new_n522_));
  INV_X1    g321(.A(G1gat), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT14), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G1gat), .B(G8gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n521_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n520_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n531_), .B(new_n520_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT80), .ZN(new_n541_));
  XOR2_X1   g340(.A(G113gat), .B(G141gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT79), .ZN(new_n543_));
  XOR2_X1   g342(.A(G169gat), .B(G197gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n541_), .B(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n517_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n439_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n487_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(new_n532_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(KEYINPUT76), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n551_), .A2(KEYINPUT76), .ZN(new_n553_));
  XOR2_X1   g352(.A(G127gat), .B(G155gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT16), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n558_));
  OR4_X1    g357(.A1(new_n552_), .A2(new_n553_), .A3(new_n557_), .A4(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n557_), .B(KEYINPUT17), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n551_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT78), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(KEYINPUT78), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n559_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n461_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n565_), .B(new_n520_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT34), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n570_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n497_), .A2(new_n501_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n565_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n576_), .B2(new_n521_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n566_), .A2(new_n573_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n578_), .A2(KEYINPUT71), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n576_), .A2(KEYINPUT70), .A3(new_n521_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT70), .ZN(new_n581_));
  INV_X1    g380(.A(new_n521_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n581_), .B1(new_n502_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(KEYINPUT71), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n579_), .A2(new_n580_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n577_), .B1(new_n585_), .B2(new_n571_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G134gat), .B(G162gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT72), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n589_), .B(KEYINPUT36), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT73), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n594_), .B1(new_n586_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n564_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n548_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT102), .ZN(new_n601_));
  AOI21_X1  g400(.A(KEYINPUT102), .B1(new_n548_), .B2(new_n599_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n393_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G1gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n596_), .B(KEYINPUT74), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n586_), .A2(new_n607_), .ZN(new_n608_));
  AOI211_X1 g407(.A(new_n577_), .B(new_n592_), .C1(new_n585_), .C2(new_n571_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT37), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT37), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n594_), .B(new_n611_), .C1(new_n586_), .C2(new_n596_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n564_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n548_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT100), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n548_), .A2(new_n617_), .A3(new_n614_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n394_), .A2(G1gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT101), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n616_), .A2(new_n622_), .A3(new_n618_), .A4(new_n619_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(KEYINPUT38), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n606_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT38), .B1(new_n621_), .B2(new_n623_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT103), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n624_), .A4(new_n606_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(G1324gat));
  NAND4_X1  g430(.A1(new_n616_), .A2(new_n522_), .A3(new_n294_), .A4(new_n618_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n600_), .A2(new_n294_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n633_), .A2(new_n634_), .A3(G8gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n633_), .B2(G8gat), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n637_), .B(new_n638_), .Z(G1325gat));
  INV_X1    g438(.A(new_n615_), .ZN(new_n640_));
  INV_X1    g439(.A(G15gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n368_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n604_), .B2(new_n368_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(KEYINPUT41), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(KEYINPUT41), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(G1326gat));
  INV_X1    g445(.A(G22gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n423_), .B(KEYINPUT105), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n640_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n648_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(new_n647_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n652_), .A2(KEYINPUT42), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(KEYINPUT42), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n650_), .B1(new_n653_), .B2(new_n654_), .ZN(G1327gat));
  INV_X1    g454(.A(new_n564_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n597_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n548_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G29gat), .B1(new_n658_), .B2(new_n393_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n353_), .A2(new_n294_), .A3(new_n393_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n434_), .B1(new_n433_), .B2(new_n353_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n368_), .B1(new_n662_), .B2(new_n435_), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT43), .B(new_n613_), .C1(new_n663_), .C2(new_n396_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n610_), .A2(new_n612_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n439_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n547_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n664_), .A2(new_n667_), .A3(new_n668_), .A4(new_n564_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n664_), .A2(new_n667_), .A3(new_n564_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(KEYINPUT44), .A4(new_n668_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT106), .B1(new_n669_), .B2(new_n670_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n393_), .A2(G29gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n659_), .B1(new_n676_), .B2(new_n677_), .ZN(G1328gat));
  NOR2_X1   g477(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n679_));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n676_), .B2(new_n294_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n658_), .A2(new_n680_), .A3(new_n294_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n679_), .B1(new_n681_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n679_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n684_), .ZN(new_n687_));
  AOI221_X4 g486(.A(new_n295_), .B1(new_n670_), .B2(new_n669_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n686_), .B(new_n687_), .C1(new_n688_), .C2(new_n680_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n685_), .A2(new_n689_), .ZN(G1329gat));
  NAND2_X1  g489(.A1(new_n368_), .A2(G43gat), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n691_), .B(new_n671_), .C1(new_n675_), .C2(new_n674_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G43gat), .B1(new_n658_), .B2(new_n368_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT47), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n691_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n676_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT47), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n698_), .ZN(G1330gat));
  AOI21_X1  g498(.A(G50gat), .B1(new_n658_), .B2(new_n649_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n423_), .A2(G50gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n676_), .B2(new_n701_), .ZN(G1331gat));
  NOR2_X1   g501(.A1(new_n439_), .A2(new_n546_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(KEYINPUT109), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(new_n517_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(KEYINPUT109), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n614_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(G57gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n393_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n599_), .A2(new_n516_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n439_), .A2(new_n546_), .A3(new_n712_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n713_), .A2(KEYINPUT110), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(KEYINPUT110), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(new_n393_), .A3(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n716_), .B2(new_n710_), .ZN(G1332gat));
  NAND3_X1  g516(.A1(new_n714_), .A2(new_n715_), .A3(new_n294_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(G64gat), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G64gat), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n295_), .A2(G64gat), .ZN(new_n722_));
  OAI22_X1  g521(.A1(new_n720_), .A2(new_n721_), .B1(new_n708_), .B2(new_n722_), .ZN(G1333gat));
  NAND3_X1  g522(.A1(new_n709_), .A2(new_n356_), .A3(new_n368_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT49), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n714_), .A2(new_n715_), .A3(new_n368_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(G71gat), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n725_), .A3(G71gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(G1334gat));
  NAND3_X1  g528(.A1(new_n714_), .A2(new_n715_), .A3(new_n649_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(G78gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n730_), .B2(G78gat), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n648_), .A2(G78gat), .ZN(new_n734_));
  OAI22_X1  g533(.A1(new_n732_), .A2(new_n733_), .B1(new_n708_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI221_X1 g536(.A(KEYINPUT112), .B1(new_n708_), .B2(new_n734_), .C1(new_n733_), .C2(new_n732_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1335gat));
  NOR2_X1   g538(.A1(new_n517_), .A2(new_n546_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n664_), .A2(new_n667_), .A3(new_n564_), .A4(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n394_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n707_), .A2(new_n657_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n393_), .A2(new_n455_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n742_), .B1(new_n743_), .B2(new_n744_), .ZN(G1336gat));
  OAI21_X1  g544(.A(G92gat), .B1(new_n741_), .B2(new_n295_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n294_), .A2(new_n456_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n743_), .B2(new_n747_), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n741_), .B2(new_n438_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n446_), .A2(new_n448_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n368_), .A2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n743_), .B2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g552(.A(G106gat), .B1(new_n741_), .B2(new_n353_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(KEYINPUT113), .A3(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n353_), .A2(G106gat), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n705_), .A2(new_n657_), .A3(new_n706_), .A4(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT52), .B1(new_n754_), .B2(KEYINPUT113), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n754_), .A2(KEYINPUT113), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n760_), .B(new_n761_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n762_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT53), .B1(new_n765_), .B2(new_n759_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  INV_X1    g566(.A(G113gat), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n516_), .A2(new_n546_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n614_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n614_), .B2(new_n770_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n502_), .A2(new_n503_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n440_), .A2(new_n319_), .A3(KEYINPUT114), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n774_), .A2(new_n488_), .A3(new_n493_), .A4(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n504_), .B2(new_n775_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n504_), .A2(new_n441_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n509_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n509_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n781_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n509_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n534_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n537_), .A2(new_n538_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  MUX2_X1   g591(.A(new_n792_), .B(new_n540_), .S(new_n545_), .Z(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n510_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT58), .B1(new_n789_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT116), .B1(new_n796_), .B2(new_n666_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n509_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n783_), .B2(new_n782_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n794_), .B1(new_n800_), .B2(new_n788_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n798_), .B(new_n613_), .C1(new_n801_), .C2(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(KEYINPUT58), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n797_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n546_), .A2(new_n510_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n787_), .B2(new_n782_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n512_), .A2(new_n793_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n597_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n809_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n804_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n773_), .B1(new_n813_), .B2(new_n564_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n354_), .A2(new_n438_), .A3(new_n394_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT117), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n546_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n768_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n820_), .A2(KEYINPUT118), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n817_), .A2(KEYINPUT119), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n816_), .A2(new_n823_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n822_), .A2(new_n824_), .A3(KEYINPUT59), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n804_), .A2(new_n812_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n810_), .B1(new_n826_), .B2(KEYINPUT120), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n804_), .A2(new_n828_), .A3(new_n812_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n656_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n825_), .B1(new_n830_), .B2(new_n773_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT59), .B1(new_n814_), .B2(new_n817_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n831_), .A2(G113gat), .A3(new_n546_), .A4(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n820_), .A2(KEYINPUT118), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n821_), .A2(new_n833_), .A3(new_n834_), .ZN(G1340gat));
  NAND2_X1  g634(.A1(new_n826_), .A2(KEYINPUT120), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(new_n811_), .A3(new_n829_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n773_), .B1(new_n837_), .B2(new_n564_), .ZN(new_n838_));
  OR3_X1    g637(.A1(new_n822_), .A2(KEYINPUT59), .A3(new_n824_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n516_), .B(new_n832_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n831_), .A2(KEYINPUT122), .A3(new_n516_), .A4(new_n832_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(G120gat), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n818_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT60), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT121), .B1(new_n846_), .B2(G120gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(G120gat), .B1(new_n516_), .B2(new_n846_), .ZN(new_n848_));
  MUX2_X1   g647(.A(new_n847_), .B(KEYINPUT121), .S(new_n848_), .Z(new_n849_));
  NAND2_X1  g648(.A1(new_n845_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n844_), .A2(new_n850_), .ZN(G1341gat));
  INV_X1    g650(.A(G127gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n564_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n831_), .A2(new_n832_), .A3(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n818_), .B2(new_n564_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n854_), .A2(KEYINPUT123), .A3(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1342gat));
  NAND3_X1  g659(.A1(new_n831_), .A2(new_n613_), .A3(new_n832_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G134gat), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n597_), .A2(G134gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n818_), .B2(new_n863_), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n814_), .A2(new_n368_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n353_), .A2(new_n294_), .A3(new_n394_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n819_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n297_), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n517_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n298_), .ZN(G1345gat));
  OAI21_X1  g670(.A(KEYINPUT124), .B1(new_n867_), .B2(new_n564_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n865_), .A2(new_n873_), .A3(new_n656_), .A4(new_n866_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n872_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1346gat));
  OAI21_X1  g677(.A(G162gat), .B1(new_n867_), .B2(new_n666_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n597_), .A2(G162gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n867_), .B2(new_n880_), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n838_), .A2(new_n649_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n295_), .A2(new_n395_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT22), .B(G169gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n546_), .A2(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT125), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n882_), .A2(new_n883_), .A3(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n648_), .B(new_n883_), .C1(new_n830_), .C2(new_n773_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n888_), .B(G169gat), .C1(new_n889_), .C2(new_n819_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n773_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n804_), .A2(new_n828_), .A3(new_n812_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n828_), .B1(new_n804_), .B2(new_n812_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n893_), .A2(new_n894_), .A3(new_n810_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n892_), .B1(new_n895_), .B2(new_n656_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n896_), .A2(new_n546_), .A3(new_n648_), .A4(new_n883_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n888_), .B1(new_n897_), .B2(G169gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n887_), .B1(new_n891_), .B2(new_n898_), .ZN(G1348gat));
  NOR2_X1   g698(.A1(new_n814_), .A2(new_n423_), .ZN(new_n900_));
  AND4_X1   g699(.A1(G176gat), .A2(new_n900_), .A3(new_n516_), .A4(new_n883_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n882_), .A2(new_n516_), .A3(new_n883_), .ZN(new_n902_));
  INV_X1    g701(.A(G176gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1349gat));
  NAND2_X1  g703(.A1(new_n656_), .A2(new_n883_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G183gat), .B1(new_n900_), .B2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n212_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n882_), .B2(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n889_), .B2(new_n666_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n598_), .A2(new_n213_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n889_), .B2(new_n911_), .ZN(G1351gat));
  NOR3_X1   g711(.A1(new_n295_), .A2(new_n353_), .A3(new_n393_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n814_), .A2(new_n368_), .A3(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n546_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n516_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g718(.A(KEYINPUT63), .B(G211gat), .Z(new_n920_));
  NAND3_X1  g719(.A1(new_n915_), .A2(new_n656_), .A3(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n921_), .A2(new_n922_), .ZN(new_n924_));
  AOI211_X1 g723(.A(KEYINPUT63), .B(G211gat), .C1(new_n915_), .C2(new_n656_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(G1354gat));
  NAND3_X1  g725(.A1(new_n915_), .A2(new_n222_), .A3(new_n598_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n915_), .A2(new_n613_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n928_), .B2(new_n222_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT127), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n927_), .B(new_n931_), .C1(new_n928_), .C2(new_n222_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1355gat));
endmodule


