//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G190gat), .B(G218gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G29gat), .B(G36gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n212_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(new_n210_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n220_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NOR4_X1   g023(.A1(new_n221_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n219_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  AND3_X1   g025(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n222_), .A2(new_n220_), .A3(new_n223_), .ZN(new_n230_));
  INV_X1    g029(.A(G99gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(new_n223_), .A3(KEYINPUT68), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT7), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n230_), .A2(new_n233_), .A3(KEYINPUT69), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n226_), .A2(new_n229_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G85gat), .ZN(new_n236_));
  INV_X1    g035(.A(G92gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G85gat), .A2(G92gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n235_), .A2(KEYINPUT8), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT9), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT9), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n239_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n238_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT67), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n231_), .A2(KEYINPUT10), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G99gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n249_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n252_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n223_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n244_), .A2(new_n256_), .A3(new_n238_), .A4(new_n246_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n248_), .A2(new_n255_), .A3(new_n229_), .A4(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n230_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n240_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT8), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n218_), .B1(new_n241_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT74), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n235_), .A2(KEYINPUT8), .A3(new_n240_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(new_n262_), .A3(new_n258_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT74), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n218_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n209_), .B1(new_n270_), .B2(KEYINPUT75), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G232gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT34), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n267_), .A2(new_n216_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n273_), .A2(new_n208_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n271_), .A2(new_n273_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n267_), .A2(new_n268_), .A3(new_n218_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n268_), .B1(new_n267_), .B2(new_n218_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT75), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  AND4_X1   g079(.A1(new_n275_), .A2(new_n280_), .A3(new_n208_), .A4(new_n273_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n202_), .B(new_n207_), .C1(new_n277_), .C2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n208_), .A3(new_n273_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n275_), .A2(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n207_), .A2(new_n202_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n207_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT36), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n275_), .A2(new_n280_), .A3(new_n208_), .A4(new_n273_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n285_), .A2(new_n286_), .A3(new_n288_), .A4(new_n289_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n282_), .A2(KEYINPUT37), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT37), .B1(new_n282_), .B2(new_n290_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G127gat), .B(G155gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(G211gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT16), .B(G183gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT17), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT78), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G15gat), .B(G22gat), .ZN(new_n301_));
  INV_X1    g100(.A(G1gat), .ZN(new_n302_));
  INV_X1    g101(.A(G8gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT14), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G1gat), .B(G8gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G231gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G71gat), .B(G78gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G57gat), .A2(G64gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT11), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G57gat), .A2(G64gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT11), .B1(new_n317_), .B2(new_n312_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n311_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n310_), .B(KEYINPUT11), .C1(new_n312_), .C2(new_n317_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n319_), .A2(new_n320_), .A3(KEYINPUT70), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT70), .B1(new_n319_), .B2(new_n320_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n309_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n300_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n319_), .A2(new_n320_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n309_), .B(new_n326_), .ZN(new_n327_));
  OR3_X1    g126(.A1(new_n327_), .A2(new_n298_), .A3(new_n297_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n293_), .A2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT79), .Z(new_n332_));
  INV_X1    g131(.A(G197gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(G204gat), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n334_), .A2(KEYINPUT93), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n333_), .A2(G204gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n336_), .B2(KEYINPUT93), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT94), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n335_), .A2(new_n337_), .B1(new_n338_), .B2(KEYINPUT21), .ZN(new_n339_));
  INV_X1    g138(.A(new_n336_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(KEYINPUT21), .A3(new_n334_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(KEYINPUT21), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n345_));
  OAI22_X1  g144(.A1(new_n339_), .A2(new_n343_), .B1(new_n345_), .B2(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT23), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n348_), .B1(new_n349_), .B2(new_n347_), .ZN(new_n350_));
  INV_X1    g149(.A(G183gat), .ZN(new_n351_));
  INV_X1    g150(.A(G190gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G169gat), .ZN(new_n356_));
  INV_X1    g155(.A(G176gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(KEYINPUT84), .A3(new_n357_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n354_), .A2(new_n355_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n349_), .A2(new_n347_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n347_), .A2(KEYINPUT23), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n368_), .B2(new_n355_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(new_n352_), .B2(KEYINPUT26), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT25), .B(G183gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT26), .B(G190gat), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n371_), .B(new_n372_), .C1(new_n373_), .C2(new_n370_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n365_), .A2(new_n369_), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n346_), .A2(new_n362_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n373_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n350_), .A2(new_n369_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n355_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n365_), .A2(new_n353_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT96), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n363_), .A2(new_n364_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n383_), .A2(KEYINPUT96), .B1(new_n357_), .B2(new_n356_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n378_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  OAI211_X1 g184(.A(KEYINPUT20), .B(new_n376_), .C1(new_n385_), .C2(new_n346_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n386_), .A2(KEYINPUT97), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT97), .B1(new_n386_), .B2(new_n390_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT100), .B(G8gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G64gat), .B(G92gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G36gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n396_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n385_), .A2(new_n346_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT98), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n346_), .B1(new_n375_), .B2(new_n362_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT98), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n385_), .A2(new_n406_), .A3(new_n346_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n402_), .A2(new_n389_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n393_), .A2(new_n400_), .A3(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n386_), .A2(new_n390_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n389_), .B1(new_n405_), .B2(new_n401_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n399_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n409_), .A2(KEYINPUT27), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT27), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n400_), .B1(new_n393_), .B2(new_n408_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n386_), .A2(new_n390_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT97), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n386_), .A2(KEYINPUT97), .A3(new_n390_), .ZN(new_n420_));
  AND4_X1   g219(.A1(new_n400_), .A2(new_n419_), .A3(new_n408_), .A4(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n415_), .B1(new_n416_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT103), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(KEYINPUT103), .B(new_n415_), .C1(new_n416_), .C2(new_n421_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n414_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT92), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT2), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(KEYINPUT92), .A2(KEYINPUT2), .ZN(new_n430_));
  OAI211_X1 g229(.A(G141gat), .B(G148gat), .C1(new_n429_), .C2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(G141gat), .ZN(new_n432_));
  INV_X1    g231(.A(G148gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n434_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n432_), .B(new_n433_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n431_), .A2(new_n439_), .A3(new_n440_), .A4(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G155gat), .B(G162gat), .Z(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n434_), .B(KEYINPUT89), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT90), .B1(new_n447_), .B2(KEYINPUT1), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT90), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT1), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(G155gat), .A4(G162gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n447_), .A2(KEYINPUT1), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G155gat), .A2(G162gat), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n446_), .B(new_n441_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n445_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G113gat), .B(G120gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G127gat), .B(G134gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G113gat), .B(G120gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(new_n459_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n461_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n456_), .A2(new_n457_), .A3(new_n462_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT101), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n460_), .B(new_n465_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT101), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n457_), .A4(new_n456_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G225gat), .A2(G233gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n456_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n466_), .A2(new_n462_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n455_), .A3(new_n445_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n477_), .A3(KEYINPUT4), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n472_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT102), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n475_), .A2(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n473_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT102), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n472_), .A2(new_n478_), .A3(new_n483_), .A4(new_n474_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(new_n236_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT0), .B(G57gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n480_), .A2(new_n482_), .A3(new_n484_), .A4(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  OR3_X1    g292(.A1(new_n456_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT28), .B1(new_n456_), .B2(KEYINPUT29), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n456_), .A2(KEYINPUT29), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(new_n346_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n494_), .B(new_n495_), .C1(new_n497_), .C2(new_n346_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G22gat), .B(G50gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G228gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G78gat), .B(G106gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n501_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G71gat), .B(G99gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G227gat), .A2(G233gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n362_), .A2(new_n512_), .A3(new_n375_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n512_), .B1(new_n362_), .B2(new_n375_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT88), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n362_), .A2(new_n375_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT30), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n513_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n516_), .A2(new_n520_), .A3(new_n469_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n469_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n511_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n516_), .A2(new_n520_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n476_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n516_), .A2(new_n520_), .A3(new_n469_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n511_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G15gat), .B(G43gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n523_), .A2(new_n528_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n531_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n508_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n531_), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n521_), .A2(new_n522_), .A3(new_n511_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n527_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n501_), .B(new_n506_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n523_), .A2(new_n528_), .A3(new_n531_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n493_), .B1(new_n534_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n400_), .A2(KEYINPUT32), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n419_), .A2(new_n408_), .A3(new_n420_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(new_n544_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n493_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT33), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n492_), .B(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(new_n399_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n472_), .A2(new_n473_), .A3(new_n478_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n481_), .A2(new_n474_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n489_), .A3(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n409_), .A2(new_n552_), .A3(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n549_), .B1(new_n551_), .B2(new_n556_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n532_), .A2(new_n533_), .A3(new_n539_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n426_), .A2(new_n542_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n332_), .A2(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n321_), .A2(new_n322_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n267_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT64), .Z(new_n566_));
  NAND4_X1  g365(.A1(new_n323_), .A2(new_n266_), .A3(new_n262_), .A4(new_n258_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n326_), .A2(new_n563_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n241_), .B2(new_n263_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n564_), .A2(new_n566_), .A3(new_n567_), .A4(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n562_), .A2(new_n567_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n566_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(G204gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT5), .B(G176gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT71), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n570_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT13), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n580_), .B(new_n581_), .C1(KEYINPUT72), .C2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT80), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n307_), .A2(new_n216_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n218_), .B2(new_n307_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n307_), .A2(new_n216_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n594_), .B1(new_n595_), .B2(new_n590_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n589_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT80), .B1(new_n591_), .B2(new_n592_), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT81), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(KEYINPUT81), .B(new_n602_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n588_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n560_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(new_n302_), .A3(new_n493_), .ZN(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n612_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT105), .ZN(new_n615_));
  AOI211_X1 g414(.A(KEYINPUT36), .B(new_n287_), .C1(new_n285_), .C2(new_n289_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n290_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n282_), .A2(KEYINPUT105), .A3(new_n290_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n559_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n608_), .A3(new_n330_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n493_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT106), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n613_), .A2(new_n614_), .A3(new_n625_), .ZN(G1324gat));
  INV_X1    g425(.A(new_n426_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n609_), .A2(new_n303_), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G8gat), .B1(new_n622_), .B2(new_n426_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT39), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n532_), .A2(new_n533_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n609_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G15gat), .B1(new_n622_), .B2(new_n638_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT41), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT108), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT108), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n640_), .A2(new_n643_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1326gat));
  INV_X1    g447(.A(G22gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n508_), .B(KEYINPUT109), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n609_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n650_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G22gat), .B1(new_n622_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT42), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(G1327gat));
  NAND2_X1  g454(.A1(new_n424_), .A2(new_n425_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n542_), .A3(new_n413_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n492_), .A2(new_n550_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n492_), .A2(new_n550_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n659_), .A2(new_n556_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n545_), .ZN(new_n662_));
  AOI211_X1 g461(.A(new_n662_), .B(new_n547_), .C1(new_n490_), .C2(new_n492_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n558_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n293_), .B1(new_n657_), .B2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n665_), .B2(KEYINPUT110), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n667_), .B(new_n668_), .C1(new_n559_), .C2(new_n293_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n588_), .A2(new_n607_), .A3(new_n330_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n666_), .A2(new_n669_), .A3(KEYINPUT44), .A4(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(new_n493_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(KEYINPUT111), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT111), .B1(new_n673_), .B2(new_n674_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT112), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT112), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(new_n672_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(G29gat), .A3(new_n681_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n282_), .A2(KEYINPUT105), .A3(new_n290_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT105), .B1(new_n282_), .B2(new_n290_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n559_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n670_), .ZN(new_n687_));
  OR3_X1    g486(.A1(new_n687_), .A2(G29gat), .A3(new_n623_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n682_), .A2(new_n688_), .ZN(G1328gat));
  INV_X1    g488(.A(new_n687_), .ZN(new_n690_));
  INV_X1    g489(.A(G36gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n627_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT45), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n671_), .A2(new_n627_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n673_), .A2(new_n674_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n694_), .B1(new_n697_), .B2(new_n675_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n693_), .B1(new_n698_), .B2(new_n691_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT113), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  OAI221_X1 g501(.A(new_n693_), .B1(new_n700_), .B2(KEYINPUT46), .C1(new_n698_), .C2(new_n691_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  INV_X1    g503(.A(G43gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n638_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n671_), .B(new_n706_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n687_), .B2(new_n638_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT47), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n707_), .A2(new_n711_), .A3(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1330gat));
  AOI21_X1  g512(.A(G50gat), .B1(new_n690_), .B2(new_n650_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n671_), .A2(G50gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n697_), .B2(new_n675_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n716_), .B2(new_n539_), .ZN(G1331gat));
  INV_X1    g516(.A(new_n588_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(new_n606_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n621_), .A2(new_n330_), .A3(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(G57gat), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n623_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n560_), .A2(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n493_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(new_n721_), .ZN(G1332gat));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(new_n726_), .A3(new_n627_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G64gat), .B1(new_n720_), .B2(new_n426_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT48), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n723_), .A2(new_n731_), .A3(new_n639_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G71gat), .B1(new_n720_), .B2(new_n638_), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n723_), .A2(new_n737_), .A3(new_n650_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G78gat), .B1(new_n720_), .B2(new_n652_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT50), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1335gat));
  NOR3_X1   g540(.A1(new_n718_), .A2(new_n606_), .A3(new_n330_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n686_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n493_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n666_), .A2(new_n669_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n742_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n493_), .A2(G85gat), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT115), .Z(new_n749_));
  AOI21_X1  g548(.A(new_n744_), .B1(new_n747_), .B2(new_n749_), .ZN(G1336gat));
  AOI21_X1  g549(.A(G92gat), .B1(new_n743_), .B2(new_n627_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n426_), .A2(new_n237_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n747_), .B2(new_n752_), .ZN(G1337gat));
  OAI21_X1  g552(.A(G99gat), .B1(new_n746_), .B2(new_n638_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n253_), .A2(new_n254_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n743_), .A2(new_n755_), .A3(new_n639_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n757_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n754_), .B(KEYINPUT117), .C1(new_n758_), .C2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g560(.A1(new_n743_), .A2(new_n223_), .A3(new_n539_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n666_), .A2(new_n669_), .A3(new_n539_), .A4(new_n742_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G106gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G106gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g567(.A(new_n606_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n293_), .A2(KEYINPUT118), .A3(new_n330_), .A4(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT37), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n282_), .A2(KEYINPUT37), .A3(new_n290_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n330_), .A4(new_n769_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n770_), .A2(new_n776_), .A3(KEYINPUT54), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n774_), .A2(new_n775_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n591_), .A2(new_n592_), .ZN(new_n781_));
  OR3_X1    g580(.A1(new_n595_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n603_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n597_), .A2(new_n598_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n603_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n582_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n569_), .A2(new_n567_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT12), .B1(new_n267_), .B2(new_n561_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n572_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT55), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n572_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n570_), .A2(KEYINPUT119), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n792_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n579_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n579_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n581_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n787_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT120), .B1(new_n804_), .B2(new_n620_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT57), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n801_), .A2(new_n581_), .A3(new_n785_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n293_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n801_), .A2(KEYINPUT58), .A3(new_n581_), .A4(new_n785_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n606_), .A2(new_n581_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n618_), .B(new_n619_), .C1(new_n814_), .C2(new_n787_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(KEYINPUT120), .A3(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n806_), .A2(new_n812_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n780_), .B1(new_n329_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n426_), .A2(new_n493_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n819_), .A2(new_n534_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821_), .B2(new_n606_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n329_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n780_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n820_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n825_), .A2(new_n639_), .A3(new_n508_), .A4(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n830_));
  NAND2_X1  g629(.A1(new_n821_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n607_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n822_), .B1(new_n832_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n718_), .B2(KEYINPUT60), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n821_), .B(new_n835_), .C1(KEYINPUT60), .C2(new_n834_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n718_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n834_), .ZN(G1341gat));
  AOI21_X1  g637(.A(G127gat), .B1(new_n821_), .B2(new_n330_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n329_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g640(.A(G134gat), .B1(new_n821_), .B2(new_n620_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n293_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845_));
  INV_X1    g644(.A(new_n541_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n826_), .A2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT122), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n819_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n847_), .B(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n579_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n579_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n803_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n786_), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n852_), .B(KEYINPUT57), .C1(new_n685_), .C2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n816_), .B1(new_n815_), .B2(KEYINPUT120), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n330_), .B1(new_n859_), .B2(new_n812_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT123), .B(new_n851_), .C1(new_n860_), .C2(new_n780_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n849_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n606_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n588_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n330_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  INV_X1    g668(.A(G162gat), .ZN(new_n870_));
  AOI211_X1 g669(.A(new_n870_), .B(new_n293_), .C1(new_n849_), .C2(new_n861_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT123), .B1(new_n825_), .B2(new_n851_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n819_), .A2(new_n845_), .A3(new_n848_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n620_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(KEYINPUT124), .A3(new_n870_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n685_), .B1(new_n849_), .B2(new_n861_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(G162gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n871_), .B1(new_n875_), .B2(new_n878_), .ZN(G1347gat));
  NOR2_X1   g678(.A1(new_n426_), .A2(new_n493_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n639_), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n819_), .A2(new_n607_), .A3(new_n650_), .A4(new_n881_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n882_), .A2(new_n356_), .ZN(new_n883_));
  INV_X1    g682(.A(G169gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT62), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1348gat));
  NOR3_X1   g688(.A1(new_n819_), .A2(new_n650_), .A3(new_n881_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G176gat), .B1(new_n890_), .B2(new_n588_), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n819_), .A2(new_n493_), .A3(new_n426_), .A4(new_n534_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n718_), .A2(new_n357_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(G1349gat));
  AOI21_X1  g693(.A(G183gat), .B1(new_n892_), .B2(new_n330_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n329_), .A2(new_n372_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n890_), .B2(new_n896_), .ZN(G1350gat));
  NAND3_X1  g696(.A1(new_n890_), .A2(new_n373_), .A3(new_n620_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n890_), .A2(new_n810_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n352_), .ZN(G1351gat));
  NAND4_X1  g699(.A1(new_n825_), .A2(new_n606_), .A3(new_n846_), .A4(new_n880_), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n901_), .A2(KEYINPUT125), .A3(new_n333_), .ZN(new_n902_));
  AOI21_X1  g701(.A(KEYINPUT125), .B1(new_n901_), .B2(new_n333_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n333_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(G1352gat));
  AND3_X1   g704(.A1(new_n825_), .A2(new_n846_), .A3(new_n880_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n588_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g707(.A(new_n329_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n909_), .B(KEYINPUT126), .Z(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n825_), .A2(new_n846_), .A3(new_n880_), .A4(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n912_), .A2(KEYINPUT127), .A3(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(KEYINPUT127), .B1(new_n912_), .B2(new_n913_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n912_), .A2(new_n913_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(G1354gat));
  AOI21_X1  g716(.A(G218gat), .B1(new_n906_), .B2(new_n620_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n810_), .A2(G218gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n906_), .B2(new_n919_), .ZN(G1355gat));
endmodule


