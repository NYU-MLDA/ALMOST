//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n824_, new_n825_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT10), .B(G99gat), .Z(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(G92gat), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT6), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n208_), .A2(new_n211_), .A3(new_n215_), .A4(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(KEYINPUT65), .B2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT7), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n217_), .B(new_n221_), .C1(new_n219_), .C2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n207_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n224_), .B1(new_n223_), .B2(new_n207_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n218_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G29gat), .B(G36gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G43gat), .B(G50gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(KEYINPUT67), .B(new_n218_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n230_), .B(new_n237_), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n232_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G232gat), .A2(G233gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(KEYINPUT34), .Z(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n238_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n247_));
  NOR4_X1   g046(.A1(new_n247_), .A2(KEYINPUT70), .A3(new_n232_), .A4(new_n245_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT35), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n246_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n244_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n250_), .B1(new_n253_), .B2(new_n248_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n206_), .B1(new_n255_), .B2(KEYINPUT71), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n257_));
  INV_X1    g056(.A(new_n206_), .ZN(new_n258_));
  AOI211_X1 g057(.A(new_n257_), .B(new_n258_), .C1(new_n252_), .C2(new_n254_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n252_), .A2(new_n254_), .A3(KEYINPUT36), .A4(new_n205_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n262_), .A2(KEYINPUT37), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(KEYINPUT37), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n260_), .A2(new_n261_), .A3(new_n263_), .A4(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n261_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(new_n262_), .A3(KEYINPUT37), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G1gat), .ZN(new_n269_));
  INV_X1    g068(.A(G8gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT14), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G15gat), .B(G22gat), .ZN(new_n274_));
  OAI211_X1 g073(.A(KEYINPUT73), .B(KEYINPUT14), .C1(new_n269_), .C2(new_n270_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G1gat), .B(G8gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G231gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G57gat), .B(G64gat), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n281_), .A2(KEYINPUT11), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(KEYINPUT11), .ZN(new_n283_));
  XOR2_X1   g082(.A(G71gat), .B(G78gat), .Z(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n283_), .A2(new_n284_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n280_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G127gat), .B(G155gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(G211gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT16), .B(G183gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n293_), .B2(KEYINPUT17), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n288_), .B(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n293_), .A2(KEYINPUT17), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n268_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT74), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G120gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT84), .B(G113gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT88), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT88), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n306_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT1), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT87), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT86), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT93), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n317_), .B(KEYINPUT3), .Z(new_n321_));
  XOR2_X1   g120(.A(new_n316_), .B(KEYINPUT2), .Z(new_n322_));
  OAI211_X1 g121(.A(new_n314_), .B(new_n311_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n305_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G225gat), .A2(G233gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n305_), .A2(new_n324_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT4), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n319_), .A2(new_n323_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n331_), .A2(new_n329_), .A3(new_n304_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n328_), .B1(new_n333_), .B2(new_n326_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G57gat), .B(G85gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G1gat), .B(G29gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n334_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G64gat), .B(G92gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT24), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT23), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354_));
  OAI211_X1 g153(.A(KEYINPUT24), .B(new_n354_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT25), .B(G183gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT26), .B(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n355_), .A2(KEYINPUT80), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT80), .B1(new_n355_), .B2(new_n358_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n351_), .B(new_n353_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n354_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT22), .B(G169gat), .ZN(new_n363_));
  INV_X1    g162(.A(G176gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n366_), .ZN(new_n368_));
  OR2_X1    g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n353_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n353_), .A2(KEYINPUT82), .A3(new_n369_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n367_), .A2(new_n368_), .A3(new_n372_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n361_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n361_), .A2(new_n374_), .A3(KEYINPUT83), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G211gat), .B(G218gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT90), .ZN(new_n380_));
  INV_X1    g179(.A(G197gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G204gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT89), .B(G204gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n383_), .B2(new_n381_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT21), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G197gat), .A2(G204gat), .ZN(new_n387_));
  OAI211_X1 g186(.A(KEYINPUT21), .B(new_n387_), .C1(new_n383_), .C2(G197gat), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n380_), .B(new_n388_), .C1(KEYINPUT21), .C2(new_n384_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n377_), .A2(new_n378_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT19), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT20), .ZN(new_n395_));
  OR3_X1    g194(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n355_), .A2(new_n358_), .A3(new_n396_), .A4(new_n353_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n370_), .A2(new_n365_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n395_), .B1(new_n390_), .B2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n392_), .A2(new_n394_), .A3(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n361_), .A2(KEYINPUT83), .A3(new_n374_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT83), .B1(new_n361_), .B2(new_n374_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n390_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT20), .B1(new_n390_), .B2(new_n399_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n394_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n347_), .B1(new_n401_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n394_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n392_), .A2(new_n409_), .A3(new_n400_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n341_), .B(new_n408_), .C1(new_n412_), .C2(new_n347_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n340_), .B1(new_n333_), .B2(new_n326_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n325_), .A2(new_n327_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(G225gat), .A3(G233gat), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n414_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n418_), .A2(new_n419_), .B1(new_n334_), .B2(new_n340_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n346_), .B1(new_n401_), .B2(new_n407_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n391_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n409_), .B1(new_n422_), .B2(new_n405_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n392_), .A2(new_n394_), .A3(new_n400_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n346_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n334_), .A2(new_n340_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n421_), .B(new_n426_), .C1(new_n427_), .C2(new_n414_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n413_), .B1(new_n420_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G15gat), .B(G43gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G71gat), .B(G99gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT30), .B1(new_n402_), .B2(new_n403_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT30), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n377_), .A2(new_n436_), .A3(new_n378_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n437_), .A3(new_n434_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n432_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n442_), .A2(new_n438_), .A3(new_n431_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n430_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n439_), .A2(new_n432_), .A3(new_n440_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n431_), .B1(new_n442_), .B2(new_n438_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(G227gat), .A4(G233gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n447_), .A3(KEYINPUT85), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n304_), .B(KEYINPUT31), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n444_), .A2(new_n447_), .A3(KEYINPUT85), .A4(new_n449_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n391_), .B1(KEYINPUT29), .B2(new_n331_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G228gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(G50gat), .B1(new_n331_), .B2(KEYINPUT29), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n458_));
  INV_X1    g257(.A(G50gat), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n319_), .A2(new_n458_), .A3(new_n459_), .A4(new_n323_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT28), .B(G22gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n457_), .A2(new_n462_), .A3(new_n460_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G78gat), .B(G106gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n457_), .A2(new_n462_), .A3(new_n460_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n462_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n456_), .B(new_n468_), .C1(new_n472_), .C2(new_n467_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n464_), .A2(KEYINPUT91), .A3(new_n465_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n466_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n456_), .B1(new_n476_), .B2(new_n468_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n429_), .A2(new_n453_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n451_), .A2(new_n452_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n425_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n421_), .A2(new_n483_), .A3(KEYINPUT27), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT27), .B1(new_n421_), .B2(new_n426_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT96), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT27), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n425_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT96), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n421_), .A2(new_n483_), .A3(KEYINPUT27), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n486_), .A2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT97), .B1(new_n494_), .B2(new_n479_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n496_));
  AOI211_X1 g295(.A(new_n496_), .B(new_n478_), .C1(new_n486_), .C2(new_n493_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n482_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n453_), .A2(new_n478_), .A3(new_n490_), .A4(new_n492_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n341_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n481_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n300_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n287_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n236_), .A2(KEYINPUT12), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G230gat), .A2(G233gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n227_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n287_), .B(KEYINPUT66), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT12), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n505_), .A2(new_n506_), .A3(new_n509_), .A4(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n509_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n507_), .A2(new_n508_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n512_), .B1(new_n506_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT68), .B(G204gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT5), .B(G176gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G120gat), .B(G148gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n516_), .A2(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT13), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(KEYINPUT13), .A3(new_n524_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(new_n381_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT76), .B(G169gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  OR3_X1    g333(.A1(new_n278_), .A2(KEYINPUT75), .A3(new_n231_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT75), .B1(new_n278_), .B2(new_n231_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n278_), .A2(new_n231_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n239_), .A2(new_n278_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n537_), .A2(new_n543_), .A3(new_n540_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n534_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n544_), .A3(new_n534_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT77), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT78), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n549_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n546_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n548_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT78), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(new_n545_), .A3(new_n550_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n530_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n503_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(new_n269_), .A3(new_n341_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT38), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n266_), .A2(KEYINPUT99), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT99), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n565_), .B(new_n261_), .C1(new_n256_), .C2(new_n259_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n502_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n559_), .A2(new_n297_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT98), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n570_), .A2(KEYINPUT98), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n569_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(G1gat), .B1(new_n573_), .B2(new_n501_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT100), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n563_), .A2(new_n575_), .ZN(G1324gat));
  INV_X1    g375(.A(new_n494_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n561_), .A2(new_n270_), .A3(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n573_), .A2(new_n494_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT39), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n579_), .A2(new_n580_), .A3(G8gat), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n579_), .B2(G8gat), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n578_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT40), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(KEYINPUT40), .B(new_n578_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(G1325gat));
  OAI21_X1  g386(.A(G15gat), .B1(new_n573_), .B2(new_n453_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT41), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n560_), .A2(G15gat), .A3(new_n453_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(G1326gat));
  OAI21_X1  g390(.A(G22gat), .B1(new_n573_), .B2(new_n479_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT42), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n479_), .A2(G22gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT101), .Z(new_n595_));
  OAI21_X1  g394(.A(new_n593_), .B1(new_n560_), .B2(new_n595_), .ZN(G1327gat));
  NAND2_X1  g395(.A1(new_n559_), .A2(new_n298_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n502_), .A2(new_n567_), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(G29gat), .B1(new_n598_), .B2(new_n341_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT44), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n265_), .A2(new_n267_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT43), .B1(new_n502_), .B2(new_n601_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n491_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n479_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n496_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n494_), .A2(KEYINPUT97), .A3(new_n479_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n453_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n490_), .A2(new_n492_), .ZN(new_n609_));
  AOI211_X1 g408(.A(new_n609_), .B(new_n479_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n501_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n480_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n268_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n597_), .B1(new_n602_), .B2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n600_), .B1(new_n615_), .B2(KEYINPUT102), .ZN(new_n616_));
  INV_X1    g415(.A(new_n597_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n613_), .B1(new_n612_), .B2(new_n268_), .ZN(new_n618_));
  AOI211_X1 g417(.A(KEYINPUT43), .B(new_n601_), .C1(new_n611_), .C2(new_n480_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n621_), .A3(KEYINPUT44), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n501_), .B1(new_n616_), .B2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n599_), .B1(new_n623_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g423(.A(G36gat), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n577_), .A2(KEYINPUT103), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n577_), .A2(KEYINPUT103), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n598_), .A2(new_n625_), .A3(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n494_), .B1(new_n616_), .B2(new_n622_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n633_), .B2(new_n625_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT46), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(KEYINPUT46), .B(new_n632_), .C1(new_n633_), .C2(new_n625_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1329gat));
  INV_X1    g437(.A(G43gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n616_), .A2(new_n622_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n640_), .B2(new_n482_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n598_), .A2(new_n639_), .A3(new_n482_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT47), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT47), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n453_), .B1(new_n616_), .B2(new_n622_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n645_), .B(new_n642_), .C1(new_n646_), .C2(new_n639_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n644_), .A2(new_n647_), .ZN(G1330gat));
  NAND3_X1  g447(.A1(new_n598_), .A2(new_n459_), .A3(new_n478_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n640_), .A2(new_n478_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n650_), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT105), .B1(new_n650_), .B2(G50gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n649_), .B1(new_n651_), .B2(new_n652_), .ZN(G1331gat));
  NOR2_X1   g452(.A1(new_n529_), .A2(new_n557_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n569_), .A2(new_n297_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(G57gat), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n501_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n503_), .A2(new_n654_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n341_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n657_), .B1(new_n660_), .B2(new_n656_), .ZN(G1332gat));
  INV_X1    g460(.A(G64gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n662_), .A3(new_n629_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT48), .ZN(new_n664_));
  INV_X1    g463(.A(new_n655_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n629_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n664_), .B1(new_n666_), .B2(G64gat), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT48), .B(new_n662_), .C1(new_n665_), .C2(new_n629_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n663_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT106), .ZN(G1333gat));
  OAI21_X1  g469(.A(G71gat), .B1(new_n655_), .B2(new_n453_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT107), .B(KEYINPUT49), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n453_), .A2(G71gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n658_), .B2(new_n674_), .ZN(G1334gat));
  OAI21_X1  g474(.A(G78gat), .B1(new_n655_), .B2(new_n479_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT50), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n479_), .A2(G78gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n658_), .B2(new_n678_), .ZN(G1335gat));
  NOR3_X1   g478(.A1(new_n529_), .A2(new_n557_), .A3(new_n297_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n612_), .A2(new_n568_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G85gat), .B1(new_n681_), .B2(new_n341_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n602_), .A2(new_n614_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(new_n680_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT108), .ZN(new_n685_));
  INV_X1    g484(.A(new_n214_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n501_), .B2(new_n212_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n682_), .B1(new_n685_), .B2(new_n687_), .ZN(G1336gat));
  AOI21_X1  g487(.A(G92gat), .B1(new_n681_), .B2(new_n577_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT109), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n685_), .A2(new_n629_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(G92gat), .ZN(G1337gat));
  NAND2_X1  g491(.A1(new_n684_), .A2(new_n482_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G99gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n681_), .A2(new_n209_), .A3(new_n482_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1338gat));
  NAND3_X1  g498(.A1(new_n681_), .A2(new_n210_), .A3(new_n478_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n683_), .A2(new_n478_), .A3(new_n680_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT52), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(G106gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n701_), .B2(G106gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g505(.A1(KEYINPUT117), .A2(G113gat), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT59), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n539_), .A2(new_n540_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n534_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n537_), .A2(new_n543_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n709_), .B(new_n710_), .C1(new_n540_), .C2(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(new_n547_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n523_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT113), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n523_), .A2(new_n716_), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n512_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT55), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n505_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(G230gat), .A3(G233gat), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT55), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n512_), .A2(new_n719_), .A3(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n721_), .A2(new_n723_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT56), .B1(new_n726_), .B2(new_n521_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(KEYINPUT56), .A3(new_n521_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n718_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT58), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n718_), .B(KEYINPUT58), .C1(new_n727_), .C2(new_n728_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n268_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n525_), .A2(new_n713_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n728_), .A2(new_n727_), .A3(KEYINPUT112), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n726_), .A2(new_n521_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT56), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(KEYINPUT112), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n522_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n734_), .B1(new_n735_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT57), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n567_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(new_n567_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n733_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n298_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n265_), .A2(new_n267_), .A3(new_n529_), .A4(new_n297_), .ZN(new_n747_));
  OR3_X1    g546(.A1(new_n747_), .A2(KEYINPUT54), .A3(new_n557_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT54), .B1(new_n747_), .B2(new_n557_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n498_), .A2(new_n501_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT116), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n752_), .A2(KEYINPUT116), .ZN(new_n754_));
  AND4_X1   g553(.A1(new_n708_), .A2(new_n751_), .A3(new_n753_), .A4(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT117), .B1(new_n557_), .B2(G113gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n745_), .A2(KEYINPUT114), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n733_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n298_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n750_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n752_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(KEYINPUT115), .A3(KEYINPUT59), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n764_));
  INV_X1    g563(.A(new_n752_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n760_), .B2(new_n750_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n766_), .B2(new_n708_), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n755_), .B(new_n756_), .C1(new_n763_), .C2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G113gat), .B1(new_n766_), .B2(new_n557_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n707_), .B1(new_n768_), .B2(new_n769_), .ZN(G1340gat));
  INV_X1    g569(.A(KEYINPUT60), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n529_), .B2(G120gat), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n766_), .B(new_n772_), .C1(new_n771_), .C2(G120gat), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n529_), .B(new_n755_), .C1(new_n763_), .C2(new_n767_), .ZN(new_n774_));
  INV_X1    g573(.A(G120gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(G1341gat));
  AOI21_X1  g575(.A(G127gat), .B1(new_n766_), .B2(new_n297_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n755_), .B1(new_n763_), .B2(new_n767_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n297_), .A2(G127gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n777_), .B1(new_n778_), .B2(new_n779_), .ZN(G1342gat));
  AOI21_X1  g579(.A(G134gat), .B1(new_n766_), .B2(new_n568_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n268_), .A2(G134gat), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT118), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n781_), .B1(new_n778_), .B2(new_n783_), .ZN(G1343gat));
  NOR2_X1   g583(.A1(new_n482_), .A2(new_n479_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n628_), .A2(new_n341_), .A3(new_n785_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT119), .Z(new_n787_));
  NAND2_X1  g586(.A1(new_n761_), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n788_), .A2(new_n558_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT120), .B(G141gat), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1344gat));
  NOR2_X1   g590(.A1(new_n788_), .A2(new_n529_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(G148gat), .Z(G1345gat));
  NAND3_X1  g592(.A1(new_n761_), .A2(new_n297_), .A3(new_n787_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n794_), .A2(G155gat), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(G155gat), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n796_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1346gat));
  INV_X1    g599(.A(G162gat), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n788_), .A2(new_n801_), .A3(new_n601_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n761_), .A2(new_n568_), .A3(new_n787_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(new_n803_), .ZN(G1347gat));
  NAND2_X1  g603(.A1(new_n629_), .A2(new_n501_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(new_n453_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n558_), .A2(new_n478_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n751_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT122), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT122), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n751_), .A2(new_n810_), .A3(new_n806_), .A4(new_n807_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(G169gat), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT123), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n809_), .A2(KEYINPUT123), .A3(G169gat), .A4(new_n811_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(KEYINPUT62), .A3(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n751_), .A2(new_n806_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n363_), .A3(new_n807_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n812_), .A2(new_n813_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n818_), .A3(new_n820_), .ZN(G1348gat));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n479_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G176gat), .B1(new_n823_), .B2(new_n530_), .ZN(new_n824_));
  AND4_X1   g623(.A1(G176gat), .A2(new_n761_), .A3(new_n530_), .A4(new_n479_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n806_), .B2(new_n825_), .ZN(G1349gat));
  NOR2_X1   g625(.A1(new_n822_), .A2(new_n298_), .ZN(new_n827_));
  MUX2_X1   g626(.A(G183gat), .B(new_n356_), .S(new_n827_), .Z(G1350gat));
  NAND3_X1  g627(.A1(new_n823_), .A2(new_n568_), .A3(new_n357_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G190gat), .B1(new_n822_), .B2(new_n601_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n830_), .A2(KEYINPUT124), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(KEYINPUT124), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n829_), .B1(new_n831_), .B2(new_n832_), .ZN(G1351gat));
  NAND4_X1  g632(.A1(new_n761_), .A2(new_n501_), .A3(new_n785_), .A4(new_n629_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n381_), .B1(new_n834_), .B2(new_n558_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT126), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT126), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n837_), .B(new_n381_), .C1(new_n834_), .C2(new_n558_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n785_), .ZN(new_n839_));
  AOI211_X1 g638(.A(new_n839_), .B(new_n805_), .C1(new_n760_), .C2(new_n750_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(G197gat), .A3(new_n557_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n840_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n557_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n836_), .A2(new_n838_), .B1(new_n843_), .B2(new_n844_), .ZN(G1352gat));
  NAND2_X1  g644(.A1(new_n840_), .A2(new_n530_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G204gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n383_), .B2(new_n846_), .ZN(G1353gat));
  NOR2_X1   g647(.A1(new_n834_), .A2(new_n298_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT127), .ZN(new_n850_));
  NOR2_X1   g649(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n849_), .A2(new_n850_), .A3(new_n852_), .A4(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n840_), .A2(new_n297_), .A3(new_n853_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT127), .B1(new_n855_), .B2(new_n851_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n851_), .B1(new_n834_), .B2(new_n298_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n854_), .A2(new_n856_), .A3(new_n857_), .ZN(G1354gat));
  AOI21_X1  g657(.A(G218gat), .B1(new_n840_), .B2(new_n568_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n268_), .A2(G218gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n840_), .B2(new_n860_), .ZN(G1355gat));
endmodule


