//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  INV_X1    g003(.A(G218gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G211gat), .ZN(new_n206_));
  INV_X1    g005(.A(G211gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G218gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n204_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G197gat), .A2(G204gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(G197gat), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(new_n211_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n206_), .A2(new_n208_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n211_), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(G197gat), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT88), .ZN(new_n224_));
  INV_X1    g023(.A(G197gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(G204gat), .ZN(new_n226_));
  INV_X1    g025(.A(G204gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT21), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n216_), .B1(new_n220_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G183gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT25), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G183gat), .ZN(new_n235_));
  INV_X1    g034(.A(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT26), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT26), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G190gat), .ZN(new_n239_));
  AND4_X1   g038(.A1(new_n233_), .A2(new_n235_), .A3(new_n237_), .A4(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(KEYINPUT74), .A2(G169gat), .A3(G176gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT74), .B1(G169gat), .B2(G176gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT75), .B1(new_n240_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n243_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT74), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(KEYINPUT74), .A2(G169gat), .A3(G176gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n233_), .A2(new_n235_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n237_), .A2(new_n239_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n251_), .B(new_n252_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT23), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(G183gat), .A3(G190gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT23), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n256_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n245_), .A2(new_n255_), .A3(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n241_), .A2(new_n242_), .ZN(new_n263_));
  INV_X1    g062(.A(G169gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT22), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT22), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(G169gat), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT76), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n260_), .A2(new_n258_), .A3(KEYINPUT77), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT77), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n273_), .A2(new_n257_), .A3(G183gat), .A4(G190gat), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n272_), .B(new_n274_), .C1(G183gat), .C2(G190gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT76), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n263_), .A2(new_n269_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n271_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n231_), .A2(new_n262_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n260_), .A2(new_n258_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n270_), .A2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n247_), .B1(new_n246_), .B2(new_n256_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n283_), .A2(new_n274_), .A3(new_n272_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT91), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n253_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT92), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n238_), .A2(G190gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n236_), .A2(KEYINPUT26), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n233_), .A2(new_n235_), .A3(KEYINPUT91), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n237_), .A2(new_n239_), .A3(KEYINPUT92), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n286_), .A2(new_n290_), .A3(new_n291_), .A4(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n282_), .B1(new_n284_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT20), .B1(new_n294_), .B2(new_n231_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n203_), .B1(new_n280_), .B2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G8gat), .B(G36gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT18), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G64gat), .B(G92gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n262_), .A2(new_n278_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n225_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n219_), .B1(new_n302_), .B2(new_n210_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n217_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n230_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n215_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT20), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(new_n294_), .B2(new_n231_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n203_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n296_), .A2(new_n300_), .A3(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n312_), .A2(KEYINPUT27), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n300_), .B(KEYINPUT97), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n280_), .A2(new_n295_), .A3(new_n203_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n310_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n300_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n307_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n319_));
  AND4_X1   g118(.A1(new_n286_), .A2(new_n290_), .A3(new_n291_), .A4(new_n292_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n283_), .A2(new_n274_), .A3(new_n272_), .ZN(new_n321_));
  OAI22_X1  g120(.A1(new_n320_), .A2(new_n321_), .B1(new_n270_), .B2(new_n281_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n308_), .B1(new_n322_), .B2(new_n306_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n310_), .B1(new_n323_), .B2(new_n279_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n318_), .B1(new_n319_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n312_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n313_), .A2(new_n317_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G228gat), .A2(G233gat), .ZN(new_n329_));
  INV_X1    g128(.A(G78gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT1), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G155gat), .A3(G162gat), .ZN(new_n336_));
  OR2_X1    g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  AND2_X1   g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT82), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT82), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n338_), .A2(new_n344_), .A3(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n347_));
  AND3_X1   g146(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT83), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n350_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n337_), .A2(KEYINPUT84), .A3(new_n333_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n358_));
  AND2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n332_), .B1(new_n346_), .B2(new_n363_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n364_), .A2(G106gat), .A3(new_n231_), .ZN(new_n365_));
  INV_X1    g164(.A(G106gat), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n338_), .A2(new_n344_), .A3(new_n341_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n344_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n357_), .A2(new_n361_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n355_), .B2(new_n350_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT29), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n366_), .B1(new_n372_), .B2(new_n306_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n331_), .B1(new_n365_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(G106gat), .B1(new_n364_), .B2(new_n231_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n366_), .A3(new_n306_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n331_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G22gat), .B(G50gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT86), .ZN(new_n381_));
  NOR4_X1   g180(.A1(new_n369_), .A2(new_n371_), .A3(KEYINPUT87), .A4(KEYINPUT29), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n343_), .A2(new_n345_), .B1(new_n356_), .B2(new_n362_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(new_n332_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n381_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n346_), .A2(new_n332_), .A3(new_n363_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT87), .ZN(new_n389_));
  INV_X1    g188(.A(new_n381_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n384_), .A2(new_n383_), .A3(new_n332_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n386_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n387_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n379_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n387_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n390_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n386_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n374_), .A4(new_n378_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n395_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n328_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT78), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT30), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n262_), .A2(new_n278_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409_));
  INV_X1    g208(.A(G71gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G99gat), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n408_), .A2(new_n412_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n407_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n301_), .B(new_n412_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n406_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n417_), .A3(KEYINPUT79), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT81), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G113gat), .B(G120gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G134gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G127gat), .ZN(new_n423_));
  INV_X1    g222(.A(G127gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G134gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n425_), .A3(KEYINPUT80), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT80), .B1(new_n423_), .B2(new_n425_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n421_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n423_), .A2(new_n425_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(new_n426_), .A3(new_n420_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT31), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n419_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n415_), .A2(new_n417_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT79), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n435_), .A2(KEYINPUT81), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n434_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n346_), .A2(new_n433_), .A3(new_n429_), .A4(new_n363_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G225gat), .A2(G233gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n443_), .A2(new_n444_), .A3(KEYINPUT4), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n448_), .B(new_n434_), .C1(new_n369_), .C2(new_n371_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n445_), .B(KEYINPUT93), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n446_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G1gat), .B(G29gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G57gat), .B(G85gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n446_), .B(new_n457_), .C1(new_n447_), .C2(new_n451_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n403_), .A2(new_n442_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n395_), .A2(new_n401_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n461_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n326_), .A2(new_n327_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n317_), .A2(KEYINPUT27), .A3(new_n312_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT99), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n443_), .A2(new_n444_), .A3(KEYINPUT4), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n471_), .A2(KEYINPUT33), .A3(new_n446_), .A4(new_n457_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n443_), .A2(new_n444_), .A3(new_n450_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n458_), .A3(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n325_), .A2(new_n472_), .A3(new_n312_), .A4(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT96), .ZN(new_n477_));
  XOR2_X1   g276(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n478_));
  AND3_X1   g277(.A1(new_n460_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n460_), .B2(new_n478_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n476_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT32), .B(new_n300_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n300_), .A2(KEYINPUT32), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n296_), .A2(new_n311_), .A3(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n461_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n402_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n328_), .A2(KEYINPUT99), .A3(new_n464_), .A4(new_n463_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n469_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n462_), .B1(new_n488_), .B2(new_n442_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n490_), .B(new_n491_), .Z(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT67), .B(KEYINPUT15), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G85gat), .B(G92gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT9), .ZN(new_n497_));
  XOR2_X1   g296(.A(KEYINPUT10), .B(G99gat), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n366_), .ZN(new_n499_));
  INV_X1    g298(.A(G85gat), .ZN(new_n500_));
  INV_X1    g299(.A(G92gat), .ZN(new_n501_));
  OR3_X1    g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT9), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT6), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G99gat), .A3(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n497_), .A2(new_n499_), .A3(new_n502_), .A4(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI211_X1 g311(.A(KEYINPUT8), .B(new_n495_), .C1(new_n512_), .C2(new_n507_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT7), .ZN(new_n515_));
  INV_X1    g314(.A(G99gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n516_), .A3(new_n366_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n505_), .B1(G99gat), .B2(G106gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n503_), .A2(KEYINPUT6), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n509_), .B(new_n517_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n514_), .B1(new_n520_), .B2(new_n496_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n508_), .B1(new_n513_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n494_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT66), .B(KEYINPUT34), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G232gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT35), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n520_), .A2(new_n496_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT8), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n520_), .A2(new_n514_), .A3(new_n496_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n490_), .B(new_n491_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n508_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n523_), .A2(new_n528_), .A3(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n526_), .A2(new_n527_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n538_));
  INV_X1    g337(.A(new_n536_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n523_), .A2(new_n539_), .A3(new_n528_), .A4(new_n534_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n537_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G190gat), .B(G218gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G134gat), .B(G162gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(KEYINPUT36), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n537_), .A2(new_n538_), .A3(new_n540_), .A4(new_n545_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550_));
  INV_X1    g349(.A(new_n544_), .ZN(new_n551_));
  AOI211_X1 g350(.A(new_n550_), .B(new_n551_), .C1(new_n537_), .C2(new_n540_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT37), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n549_), .B2(new_n553_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559_));
  INV_X1    g358(.A(G1gat), .ZN(new_n560_));
  INV_X1    g359(.A(G8gat), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT14), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G1gat), .B(G8gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G57gat), .B(G64gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G71gat), .B(G78gat), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(KEYINPUT11), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(KEYINPUT11), .ZN(new_n569_));
  INV_X1    g368(.A(new_n567_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n566_), .A2(KEYINPUT11), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n568_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n565_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT69), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n574_), .B(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G127gat), .B(G155gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT70), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n583_), .A3(KEYINPUT17), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n577_), .A2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n577_), .B(new_n584_), .C1(KEYINPUT17), .C2(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n558_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G113gat), .B(G141gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT72), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G169gat), .B(G197gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n565_), .B(new_n492_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n565_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n533_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n533_), .B(new_n493_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n599_), .B(new_n595_), .C1(new_n600_), .C2(new_n598_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n593_), .B1(new_n597_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n597_), .A2(new_n601_), .A3(new_n593_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n605_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT73), .B1(new_n607_), .B2(new_n602_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT13), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G120gat), .B(G148gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT5), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G176gat), .B(G204gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(KEYINPUT65), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT64), .ZN(new_n618_));
  INV_X1    g417(.A(new_n573_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT12), .B1(new_n522_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n522_), .A2(new_n619_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n573_), .B(new_n508_), .C1(new_n513_), .C2(new_n521_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n620_), .B1(new_n623_), .B2(KEYINPUT12), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n618_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT12), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n627_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n625_), .ZN(new_n629_));
  NOR4_X1   g428(.A1(new_n628_), .A2(KEYINPUT64), .A3(new_n629_), .A4(new_n620_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n623_), .A2(new_n629_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n617_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n573_), .B1(new_n532_), .B2(new_n508_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n622_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT12), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n620_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n625_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT64), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n624_), .A2(new_n618_), .A3(new_n625_), .ZN(new_n640_));
  AND4_X1   g439(.A1(new_n632_), .A2(new_n639_), .A3(new_n640_), .A4(new_n617_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n611_), .B1(new_n633_), .B2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n631_), .A2(new_n632_), .A3(new_n617_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n639_), .A2(new_n632_), .A3(new_n640_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n617_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n646_), .A3(KEYINPUT13), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n642_), .A2(new_n647_), .ZN(new_n648_));
  NOR4_X1   g447(.A1(new_n489_), .A2(new_n589_), .A3(new_n610_), .A4(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n560_), .A3(new_n461_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT100), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n549_), .A2(new_n553_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n489_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n642_), .A2(new_n609_), .A3(new_n647_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT101), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n642_), .A2(new_n659_), .A3(new_n609_), .A4(new_n647_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n658_), .A2(new_n588_), .A3(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n656_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n560_), .B1(new_n662_), .B2(new_n461_), .ZN(new_n663_));
  OR3_X1    g462(.A1(new_n653_), .A2(new_n654_), .A3(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(new_n328_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n649_), .A2(new_n561_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n662_), .A2(new_n665_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(G8gat), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT39), .B(new_n561_), .C1(new_n662_), .C2(new_n665_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g471(.A(G15gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n442_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n649_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n662_), .A2(new_n674_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n676_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT41), .B1(new_n676_), .B2(G15gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(G1326gat));
  NOR2_X1   g478(.A1(new_n402_), .A2(G22gat), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT102), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n649_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n662_), .A2(new_n463_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(G22gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G22gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT103), .Z(G1327gat));
  NAND2_X1  g487(.A1(new_n655_), .A2(new_n587_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT106), .Z(new_n690_));
  INV_X1    g489(.A(new_n648_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n489_), .A3(new_n610_), .ZN(new_n693_));
  INV_X1    g492(.A(G29gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n461_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  INV_X1    g496(.A(new_n557_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n555_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n461_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n460_), .A2(new_n478_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT96), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n460_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n704_), .B2(new_n476_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n468_), .A2(new_n467_), .B1(new_n705_), .B2(new_n402_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n674_), .B1(new_n706_), .B2(new_n487_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n697_), .B(new_n699_), .C1(new_n707_), .C2(new_n462_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n489_), .B2(new_n558_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n658_), .A2(new_n587_), .A3(new_n660_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n658_), .A2(KEYINPUT104), .A3(new_n587_), .A4(new_n660_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n710_), .A2(new_n715_), .A3(KEYINPUT44), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT44), .B1(new_n710_), .B2(new_n715_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n461_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n696_), .B1(new_n719_), .B2(G29gat), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT105), .B(new_n694_), .C1(new_n718_), .C2(new_n461_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n695_), .B1(new_n720_), .B2(new_n721_), .ZN(G1328gat));
  XOR2_X1   g521(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n723_));
  NOR2_X1   g522(.A1(new_n328_), .A2(G36gat), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n693_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n693_), .B2(new_n724_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n716_), .A2(new_n717_), .A3(new_n328_), .ZN(new_n728_));
  INV_X1    g527(.A(G36gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n730_), .A2(new_n731_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n717_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n710_), .A2(new_n715_), .A3(KEYINPUT44), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n665_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G36gat), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n739_), .A2(new_n732_), .A3(new_n733_), .A4(new_n727_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n735_), .A2(new_n740_), .ZN(G1329gat));
  AOI21_X1  g540(.A(G43gat), .B1(new_n693_), .B2(new_n674_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n674_), .A2(G43gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n718_), .B2(new_n743_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g544(.A(G50gat), .B1(new_n693_), .B2(new_n463_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n463_), .A2(G50gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n718_), .B2(new_n747_), .ZN(G1331gat));
  NOR2_X1   g547(.A1(new_n489_), .A2(new_n609_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n589_), .A2(new_n691_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n464_), .B1(new_n751_), .B2(KEYINPUT109), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(KEYINPUT109), .B2(new_n751_), .ZN(new_n753_));
  INV_X1    g552(.A(G57gat), .ZN(new_n754_));
  AND4_X1   g553(.A1(new_n610_), .A2(new_n656_), .A3(new_n648_), .A4(new_n588_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n464_), .A2(new_n754_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n753_), .A2(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(G1332gat));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n755_), .B2(new_n665_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT48), .Z(new_n760_));
  INV_X1    g559(.A(new_n751_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n758_), .A3(new_n665_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1333gat));
  AOI21_X1  g562(.A(new_n410_), .B1(new_n755_), .B2(new_n674_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT49), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n410_), .A3(new_n674_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1334gat));
  AOI21_X1  g566(.A(new_n330_), .B1(new_n755_), .B2(new_n463_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n768_), .B(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n761_), .A2(new_n330_), .A3(new_n463_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1335gat));
  AND2_X1   g571(.A1(new_n690_), .A2(new_n648_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n749_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n500_), .B1(new_n774_), .B2(new_n464_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n691_), .A2(new_n609_), .A3(new_n588_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n710_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n461_), .A2(G85gat), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT111), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT112), .ZN(G1336gat));
  OAI21_X1  g580(.A(G92gat), .B1(new_n777_), .B2(new_n328_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n774_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n501_), .A3(new_n665_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1337gat));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n674_), .A3(new_n498_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n777_), .A2(new_n442_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n516_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g588(.A(G106gat), .B1(new_n777_), .B2(new_n402_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n790_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT52), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n402_), .A2(G106gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n773_), .A2(new_n749_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n797_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n801_));
  AND4_X1   g600(.A1(new_n792_), .A2(new_n794_), .A3(new_n800_), .A4(new_n801_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n793_), .A2(KEYINPUT52), .B1(new_n798_), .B2(new_n799_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(new_n803_), .B2(new_n792_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1339gat));
  INV_X1    g604(.A(G113gat), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n639_), .A2(new_n632_), .A3(new_n640_), .A4(new_n616_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n609_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n609_), .A2(new_n807_), .A3(KEYINPUT115), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  NOR4_X1   g611(.A1(new_n628_), .A2(new_n812_), .A3(new_n629_), .A4(new_n620_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT116), .B1(new_n624_), .B2(new_n625_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n629_), .C1(new_n628_), .C2(new_n620_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n813_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n639_), .A2(new_n812_), .A3(new_n640_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n616_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(KEYINPUT56), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n821_), .B(new_n616_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n810_), .B(new_n811_), .C1(new_n820_), .C2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n593_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(KEYINPUT117), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n599_), .A2(new_n596_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n565_), .B2(new_n494_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(KEYINPUT117), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n607_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n633_), .B2(new_n641_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n655_), .B1(new_n823_), .B2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n819_), .B(KEYINPUT56), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n830_), .A2(new_n807_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT58), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT58), .B(new_n834_), .C1(new_n820_), .C2(new_n822_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n699_), .ZN(new_n837_));
  OAI22_X1  g636(.A1(new_n832_), .A2(KEYINPUT57), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  AOI211_X1 g638(.A(new_n839_), .B(new_n655_), .C1(new_n823_), .C2(new_n831_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n587_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n691_), .A2(new_n558_), .A3(new_n610_), .A4(new_n588_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT54), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n403_), .A2(new_n442_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n461_), .A3(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n806_), .B1(new_n846_), .B2(new_n610_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT118), .B(new_n806_), .C1(new_n846_), .C2(new_n610_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n846_), .A2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n844_), .A2(KEYINPUT59), .A3(new_n461_), .A4(new_n845_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n610_), .A2(new_n806_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n849_), .A2(new_n850_), .B1(new_n854_), .B2(new_n855_), .ZN(G1340gat));
  AOI21_X1  g655(.A(new_n691_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n857_));
  INV_X1    g656(.A(G120gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n691_), .B2(KEYINPUT60), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(KEYINPUT60), .B2(new_n858_), .ZN(new_n860_));
  OAI22_X1  g659(.A1(new_n857_), .A2(new_n858_), .B1(new_n846_), .B2(new_n860_), .ZN(G1341gat));
  INV_X1    g660(.A(new_n846_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(new_n424_), .A3(new_n588_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n587_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n424_), .ZN(G1342gat));
  NAND3_X1  g664(.A1(new_n862_), .A2(new_n422_), .A3(new_n655_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n558_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n422_), .ZN(G1343gat));
  NOR3_X1   g667(.A1(new_n674_), .A2(new_n402_), .A3(new_n665_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n844_), .A2(new_n461_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n609_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n648_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n844_), .A2(new_n461_), .A3(new_n588_), .A4(new_n869_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT119), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n877_), .A2(KEYINPUT119), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n876_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n880_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n878_), .A3(new_n875_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1346gat));
  INV_X1    g683(.A(G162gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n870_), .A2(new_n885_), .A3(new_n655_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n870_), .A2(new_n699_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1347gat));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n442_), .A2(new_n461_), .A3(new_n328_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n609_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT120), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n844_), .A2(new_n892_), .A3(new_n402_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(new_n894_), .A3(G169gat), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n893_), .B2(G169gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n889_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n893_), .A2(G169gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT121), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(KEYINPUT62), .A3(new_n895_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n844_), .A2(new_n402_), .A3(new_n890_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n903_), .A2(new_n265_), .A3(new_n267_), .A4(new_n609_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n898_), .A2(new_n901_), .A3(new_n904_), .ZN(G1348gat));
  NOR2_X1   g704(.A1(new_n902_), .A2(new_n691_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n268_), .ZN(G1349gat));
  NOR2_X1   g706(.A1(new_n902_), .A2(new_n587_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(G183gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n286_), .A2(new_n291_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n908_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n902_), .B2(new_n558_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n655_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n902_), .B2(new_n913_), .ZN(G1351gat));
  NAND3_X1  g713(.A1(new_n442_), .A2(new_n464_), .A3(new_n463_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n915_), .A2(KEYINPUT122), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(KEYINPUT122), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n916_), .A2(new_n665_), .A3(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n610_), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n225_), .A2(KEYINPUT123), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n225_), .A2(KEYINPUT123), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n921_), .B2(new_n923_), .ZN(G1352gat));
  NOR2_X1   g724(.A1(new_n920_), .A2(new_n691_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n221_), .A2(new_n222_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n926_), .A2(KEYINPUT124), .A3(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G204gat), .B1(new_n920_), .B2(new_n691_), .ZN(new_n930_));
  AOI21_X1  g729(.A(KEYINPUT124), .B1(new_n926_), .B2(new_n928_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(G1353gat));
  AOI21_X1  g731(.A(new_n587_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n919_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(KEYINPUT125), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n919_), .A2(new_n936_), .A3(new_n933_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n938_), .B(new_n939_), .ZN(G1354gat));
  NAND3_X1  g739(.A1(new_n919_), .A2(G218gat), .A3(new_n699_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n942_));
  INV_X1    g741(.A(new_n918_), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n844_), .A2(new_n942_), .A3(new_n655_), .A4(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n205_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n942_), .B1(new_n919_), .B2(new_n655_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n941_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(KEYINPUT127), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n941_), .B(new_n949_), .C1(new_n945_), .C2(new_n946_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n950_), .ZN(G1355gat));
endmodule


