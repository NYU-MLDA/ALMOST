//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n958_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n970_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G197gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G204gat), .ZN(new_n207_));
  INV_X1    g006(.A(G204gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(G197gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT21), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n205_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G211gat), .B(G218gat), .Z(new_n213_));
  OAI211_X1 g012(.A(new_n213_), .B(KEYINPUT21), .C1(new_n207_), .C2(new_n209_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT1), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(new_n218_), .B2(KEYINPUT1), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT79), .ZN(new_n223_));
  INV_X1    g022(.A(G155gat), .ZN(new_n224_));
  INV_X1    g023(.A(G162gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(G155gat), .A3(G162gat), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n217_), .B1(new_n222_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G141gat), .ZN(new_n232_));
  INV_X1    g031(.A(G148gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n226_), .A2(new_n227_), .A3(new_n218_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT81), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT3), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n217_), .A2(KEYINPUT2), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT2), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n216_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n241_), .A2(new_n232_), .A3(new_n233_), .A4(KEYINPUT81), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n237_), .A2(new_n238_), .A3(new_n240_), .A4(new_n242_), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n231_), .A2(new_n234_), .B1(new_n235_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n202_), .B(new_n215_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n202_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n218_), .A2(KEYINPUT1), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT80), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT1), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n216_), .B(new_n234_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n243_), .A2(new_n235_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n245_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n212_), .A2(new_n214_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n247_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G78gat), .B(G106gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT82), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT83), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n246_), .A2(new_n257_), .A3(new_n258_), .A4(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n253_), .A2(new_n245_), .A3(new_n254_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G22gat), .B(G50gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT28), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n263_), .B(new_n265_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n246_), .A2(new_n257_), .A3(new_n261_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n260_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n269_), .B1(new_n246_), .B2(new_n257_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n270_), .B2(KEYINPUT84), .ZN(new_n271_));
  INV_X1    g070(.A(new_n261_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n253_), .A2(new_n254_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT29), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n202_), .B1(new_n274_), .B2(new_n215_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n255_), .A2(new_n247_), .A3(new_n256_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n272_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n268_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n266_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n267_), .A2(new_n271_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G71gat), .B(G99gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G176gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n286_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT75), .B(G190gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(G183gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n290_), .B(new_n291_), .C1(new_n293_), .C2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT25), .B(G183gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n300_), .B1(new_n292_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(G190gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(KEYINPUT24), .A3(new_n291_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT24), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n308_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n299_), .B1(new_n305_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT30), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n318_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(G113gat), .A2(G120gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G113gat), .A2(G120gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(G127gat), .A2(G134gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G127gat), .A2(G134gat), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT76), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n329_));
  OR2_X1    g128(.A1(G127gat), .A2(G134gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G127gat), .A2(G134gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n325_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT76), .B1(new_n326_), .B2(new_n327_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n324_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(KEYINPUT77), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n324_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n321_), .A2(new_n341_), .ZN(new_n342_));
  AOI211_X1 g141(.A(KEYINPUT77), .B(new_n324_), .C1(new_n335_), .C2(new_n334_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n334_), .A2(new_n335_), .A3(new_n324_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(new_n338_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n345_), .B2(KEYINPUT77), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n319_), .A2(new_n346_), .A3(new_n320_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G15gat), .B(G43gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT31), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n342_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n342_), .B2(new_n347_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n285_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT0), .B(G57gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G85gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(G1gat), .B(G29gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n333_), .A2(new_n336_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n254_), .A3(new_n253_), .ZN(new_n360_));
  OAI211_X1 g159(.A(KEYINPUT4), .B(new_n360_), .C1(new_n346_), .C2(new_n244_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n337_), .A2(new_n340_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n361_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n359_), .A2(new_n254_), .A3(new_n253_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n362_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n358_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n363_), .A2(new_n370_), .A3(new_n364_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n341_), .A2(new_n364_), .A3(new_n273_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n362_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT89), .B1(new_n374_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n361_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n378_), .A2(new_n372_), .A3(new_n379_), .A4(new_n358_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n373_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n342_), .A2(new_n347_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n349_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n284_), .A3(new_n351_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n354_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n308_), .A2(new_n313_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n387_), .B(new_n310_), .C1(new_n304_), .C2(new_n302_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n256_), .A2(new_n299_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT86), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(KEYINPUT24), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n312_), .A2(KEYINPUT86), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n311_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n312_), .A2(KEYINPUT86), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n390_), .A2(KEYINPUT24), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n309_), .A2(new_n394_), .A3(new_n395_), .A4(new_n291_), .ZN(new_n396_));
  INV_X1    g195(.A(G190gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT26), .ZN(new_n398_));
  AND2_X1   g197(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n303_), .B(new_n398_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n393_), .A2(new_n396_), .A3(new_n401_), .A4(new_n308_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n288_), .A2(new_n289_), .A3(KEYINPUT87), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n405_));
  OR2_X1    g204(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n406_), .B2(new_n287_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n286_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G183gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n397_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n296_), .A2(new_n297_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n291_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT88), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT87), .B1(new_n288_), .B2(new_n289_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n406_), .A2(new_n405_), .A3(new_n287_), .ZN(new_n417_));
  AOI21_X1  g216(.A(G176gat), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT88), .B1(new_n418_), .B2(new_n412_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n403_), .B1(new_n415_), .B2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(KEYINPUT20), .B(new_n389_), .C1(new_n420_), .C2(new_n256_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n422_), .B(KEYINPUT85), .Z(new_n423_));
  XOR2_X1   g222(.A(new_n423_), .B(KEYINPUT19), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n420_), .A2(new_n256_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n428_), .B1(new_n315_), .B2(new_n215_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT18), .B(G64gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(G92gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G8gat), .B(G36gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G92gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n432_), .B(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n434_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n431_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n426_), .A2(new_n430_), .A3(new_n435_), .A4(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT97), .B(KEYINPUT27), .Z(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n440_), .B(KEYINPUT95), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT93), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n402_), .B1(new_n418_), .B2(new_n412_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT92), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n402_), .B(new_n451_), .C1(new_n418_), .C2(new_n412_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n256_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n429_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n448_), .B1(new_n454_), .B2(new_n425_), .ZN(new_n455_));
  AOI211_X1 g254(.A(KEYINPUT93), .B(new_n424_), .C1(new_n453_), .C2(new_n429_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n421_), .A2(new_n425_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n447_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT96), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n442_), .A2(KEYINPUT27), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n454_), .A2(new_n425_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT93), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n454_), .A2(new_n448_), .A3(new_n425_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n458_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n446_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n442_), .A2(KEYINPUT27), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT96), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n445_), .B1(new_n462_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT99), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n443_), .A2(new_n444_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n460_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(KEYINPUT96), .A3(new_n468_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT99), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  AOI211_X1 g276(.A(new_n281_), .B(new_n386_), .C1(new_n471_), .C2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n369_), .A2(new_n479_), .A3(new_n372_), .A4(new_n358_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n380_), .A2(KEYINPUT33), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n361_), .A2(new_n362_), .A3(new_n375_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n358_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n371_), .A2(new_n376_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n441_), .A2(new_n442_), .A3(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n482_), .A2(new_n483_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n483_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n435_), .A2(new_n439_), .A3(KEYINPUT32), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n491_), .B(KEYINPUT91), .Z(new_n492_));
  NOR2_X1   g291(.A1(new_n431_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n378_), .A2(new_n372_), .A3(new_n379_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n485_), .ZN(new_n495_));
  AOI221_X4 g294(.A(new_n493_), .B1(new_n466_), .B2(new_n491_), .C1(new_n495_), .C2(new_n380_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n489_), .A2(new_n490_), .A3(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT94), .B1(new_n497_), .B2(new_n281_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n373_), .A2(new_n280_), .A3(new_n381_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n499_), .B(new_n445_), .C1(new_n462_), .C2(new_n469_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT98), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT98), .B1(new_n475_), .B2(new_n499_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n380_), .A2(KEYINPUT33), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n380_), .A2(KEYINPUT33), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n488_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT90), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n466_), .A2(new_n491_), .ZN(new_n509_));
  OAI221_X1 g308(.A(new_n509_), .B1(new_n431_), .B2(new_n492_), .C1(new_n373_), .C2(new_n381_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n482_), .A2(new_n483_), .A3(new_n488_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n280_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n498_), .A2(new_n504_), .A3(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n354_), .A2(new_n385_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n478_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G29gat), .B(G36gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G43gat), .ZN(new_n521_));
  INV_X1    g320(.A(G50gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n520_), .A2(G43gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(G43gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(G50gat), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT73), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G1gat), .A2(G8gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT14), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G1gat), .B(G8gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n528_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT69), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n527_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT15), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n527_), .B(KEYINPUT69), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT15), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n519_), .B(new_n536_), .C1(new_n543_), .C2(new_n534_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n528_), .B(new_n535_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(G229gat), .A3(G233gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G169gat), .B(G197gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT74), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G113gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(new_n232_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G71gat), .B(G78gat), .ZN(new_n560_));
  OR3_X1    g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(new_n560_), .A3(KEYINPUT11), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT6), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT65), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G85gat), .B(G92gat), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT9), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT10), .B(G99gat), .Z(new_n571_));
  INV_X1    g370(.A(G106gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n436_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n436_), .A2(KEYINPUT64), .ZN(new_n575_));
  OAI21_X1  g374(.A(G85gat), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n567_), .A2(new_n570_), .A3(new_n573_), .A4(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT7), .ZN(new_n579_));
  AOI211_X1 g378(.A(KEYINPUT8), .B(new_n568_), .C1(new_n567_), .C2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n565_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n569_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT8), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n563_), .B(new_n577_), .C1(new_n580_), .C2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT67), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT67), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(new_n589_), .A3(new_n586_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n580_), .A2(KEYINPUT66), .A3(new_n584_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT66), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT8), .B1(new_n567_), .B2(new_n579_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n569_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n595_), .B2(new_n583_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n577_), .B1(new_n592_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n563_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(KEYINPUT12), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600_));
  INV_X1    g399(.A(new_n577_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n595_), .B2(new_n583_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n600_), .B1(new_n602_), .B2(new_n563_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n591_), .A2(new_n599_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n586_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n602_), .A2(new_n563_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n585_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n605_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n208_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT5), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(new_n286_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n604_), .A2(new_n608_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n612_), .B1(new_n604_), .B2(new_n608_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n556_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(KEYINPUT68), .A3(new_n613_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT13), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n518_), .A2(new_n555_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n563_), .B(new_n534_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT17), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT16), .B(G183gat), .ZN(new_n629_));
  INV_X1    g428(.A(G211gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G127gat), .B(G155gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n627_), .B1(new_n628_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(KEYINPUT17), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n627_), .B2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT72), .Z(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT66), .B1(new_n580_), .B2(new_n584_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n595_), .A2(new_n593_), .A3(new_n583_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n601_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n602_), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n543_), .A2(new_n640_), .B1(new_n527_), .B2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT70), .B1(new_n543_), .B2(new_n640_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(G232gat), .A2(G233gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT34), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(KEYINPUT35), .A3(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(KEYINPUT35), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n642_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT71), .B(G134gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(G162gat), .ZN(new_n651_));
  XOR2_X1   g450(.A(G190gat), .B(G218gat), .Z(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT36), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n653_), .A2(new_n654_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n646_), .A2(new_n642_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n649_), .A2(new_n655_), .A3(new_n656_), .A4(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n657_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n654_), .B(new_n653_), .C1(new_n659_), .C2(new_n648_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT37), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n658_), .A2(KEYINPUT37), .A3(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n624_), .A2(new_n637_), .A3(new_n666_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n667_), .A2(G1gat), .A3(new_n382_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT38), .ZN(new_n669_));
  INV_X1    g468(.A(new_n478_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n512_), .A2(new_n513_), .A3(new_n280_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n513_), .B1(new_n512_), .B2(new_n280_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n500_), .A2(new_n501_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n475_), .A2(KEYINPUT98), .A3(new_n499_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n671_), .A2(new_n672_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n670_), .B1(new_n676_), .B2(new_n516_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n623_), .A2(new_n555_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n637_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n661_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n382_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G1gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n668_), .A2(KEYINPUT38), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n669_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1324gat));
  XOR2_X1   g488(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n667_), .ZN(new_n692_));
  INV_X1    g491(.A(G8gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n471_), .A2(new_n477_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n692_), .A2(new_n693_), .A3(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n681_), .A2(new_n680_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n624_), .A2(new_n697_), .A3(new_n695_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT39), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(G8gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G8gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n696_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT102), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n702_), .A2(KEYINPUT102), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n691_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n702_), .A2(KEYINPUT102), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(new_n690_), .A3(new_n703_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1325gat));
  INV_X1    g508(.A(G15gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n682_), .B2(new_n516_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT41), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n692_), .A2(new_n710_), .A3(new_n516_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1326gat));
  INV_X1    g513(.A(G22gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n682_), .B2(new_n281_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT42), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n692_), .A2(new_n715_), .A3(new_n281_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1327gat));
  NAND2_X1  g518(.A1(new_n681_), .A2(new_n680_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT104), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n679_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G29gat), .B1(new_n722_), .B2(new_n683_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n677_), .B2(new_n665_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n518_), .A2(KEYINPUT43), .A3(new_n666_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n678_), .A2(new_n680_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT103), .B(KEYINPUT44), .C1(new_n727_), .C2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n677_), .A2(new_n724_), .A3(new_n665_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT43), .B1(new_n518_), .B2(new_n666_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(KEYINPUT103), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(KEYINPUT103), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n382_), .B1(new_n729_), .B2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n723_), .B1(new_n736_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g536(.A(G36gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n722_), .A2(new_n738_), .A3(new_n695_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT45), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n694_), .B1(new_n729_), .B2(new_n735_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(new_n738_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n742_), .B(new_n744_), .ZN(G1329gat));
  NOR4_X1   g544(.A1(new_n679_), .A2(new_n721_), .A3(G43gat), .A4(new_n517_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n735_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n734_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n516_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n746_), .B1(new_n749_), .B2(G43gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n722_), .B2(new_n281_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n280_), .B1(new_n729_), .B2(new_n735_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(G50gat), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n621_), .A2(new_n622_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(new_n554_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n677_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n663_), .A2(new_n637_), .A3(new_n664_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G57gat), .B1(new_n759_), .B2(new_n683_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n757_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(new_n382_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n760_), .B1(new_n763_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g563(.A(G64gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n759_), .A2(new_n765_), .A3(new_n695_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G64gat), .B1(new_n762_), .B2(new_n694_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(KEYINPUT48), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(KEYINPUT48), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT106), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n766_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1333gat));
  INV_X1    g573(.A(G71gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n761_), .B2(new_n516_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT49), .Z(new_n777_));
  NAND3_X1  g576(.A1(new_n759_), .A2(new_n775_), .A3(new_n516_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n761_), .A2(new_n281_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G78gat), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(KEYINPUT107), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(KEYINPUT107), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n784_));
  OR3_X1    g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(G78gat), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n759_), .A2(new_n786_), .A3(new_n281_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n784_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n787_), .A3(new_n788_), .ZN(G1335gat));
  NOR2_X1   g588(.A1(new_n757_), .A2(new_n721_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n683_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n727_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n756_), .A2(new_n680_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT108), .B1(new_n725_), .B2(new_n726_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n793_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(new_n683_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n791_), .B1(new_n798_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g598(.A(G92gat), .B1(new_n790_), .B2(new_n695_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n436_), .A2(KEYINPUT64), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n695_), .B1(new_n575_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT109), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n800_), .B1(new_n797_), .B2(new_n803_), .ZN(G1337gat));
  NAND3_X1  g603(.A1(new_n790_), .A2(new_n571_), .A3(new_n516_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT110), .Z(new_n806_));
  NAND4_X1  g605(.A1(new_n793_), .A2(new_n516_), .A3(new_n795_), .A4(new_n796_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G99gat), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(G1338gat));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n280_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n572_), .B1(new_n813_), .B2(new_n795_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n812_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n281_), .B(new_n795_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n815_), .A3(G106gat), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n280_), .B(new_n794_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT113), .B(KEYINPUT52), .C1(new_n821_), .C2(new_n572_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n817_), .A2(KEYINPUT112), .A3(new_n815_), .A4(G106gat), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n816_), .A2(new_n820_), .A3(new_n822_), .A4(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n790_), .A2(new_n572_), .A3(new_n281_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT53), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n824_), .A2(new_n828_), .A3(new_n825_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1339gat));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n545_), .A2(new_n519_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n536_), .B1(new_n543_), .B2(new_n534_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n551_), .B(new_n832_), .C1(new_n833_), .C2(new_n519_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n552_), .A2(new_n834_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n616_), .A2(new_n835_), .A3(new_n618_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n591_), .A2(new_n599_), .A3(KEYINPUT55), .A4(new_n603_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT114), .ZN(new_n838_));
  INV_X1    g637(.A(new_n603_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n640_), .A2(new_n600_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n598_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(KEYINPUT55), .A4(new_n591_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n599_), .A2(new_n603_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n605_), .B1(new_n844_), .B2(new_n607_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n604_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n838_), .A2(new_n843_), .A3(new_n845_), .A4(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n612_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n851_), .A2(new_n554_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n614_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n836_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n831_), .B1(new_n855_), .B2(new_n681_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n848_), .A2(new_n849_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT56), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT56), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n848_), .A2(new_n859_), .A3(new_n849_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n858_), .A2(new_n613_), .A3(new_n835_), .A4(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n860_), .A2(new_n613_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n864_), .A2(KEYINPUT58), .A3(new_n835_), .A4(new_n858_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n865_), .A3(new_n665_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n851_), .A2(new_n554_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n867_), .A2(new_n614_), .A3(new_n853_), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT57), .B(new_n661_), .C1(new_n868_), .C2(new_n836_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n856_), .A2(new_n866_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n680_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n621_), .A2(new_n622_), .A3(new_n554_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT54), .B1(new_n873_), .B2(new_n758_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n666_), .A2(new_n872_), .A3(new_n875_), .A4(new_n637_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n281_), .B1(new_n871_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n695_), .A2(new_n382_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n516_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n555_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n883_), .A2(new_n884_), .A3(G113gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(G113gat), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT59), .B1(new_n878_), .B2(new_n881_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n870_), .A2(new_n680_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n281_), .A4(new_n880_), .ZN(new_n890_));
  OAI211_X1 g689(.A(G113gat), .B(new_n554_), .C1(new_n887_), .C2(new_n890_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n885_), .A2(new_n886_), .A3(new_n891_), .ZN(G1340gat));
  INV_X1    g691(.A(new_n882_), .ZN(new_n893_));
  INV_X1    g692(.A(G120gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n894_), .B1(new_n755_), .B2(KEYINPUT60), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n893_), .B(new_n895_), .C1(KEYINPUT60), .C2(new_n894_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n887_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n890_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n755_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n896_), .B1(new_n899_), .B2(new_n894_), .ZN(G1341gat));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n901_));
  OAI21_X1  g700(.A(G127gat), .B1(new_n680_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(G127gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT117), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n902_), .B(new_n904_), .C1(new_n887_), .C2(new_n890_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n882_), .B2(new_n680_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT118), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n905_), .A2(new_n909_), .A3(new_n906_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1342gat));
  AOI21_X1  g710(.A(G134gat), .B1(new_n893_), .B2(new_n681_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n666_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT119), .B(G134gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1343gat));
  NOR3_X1   g714(.A1(new_n888_), .A2(new_n516_), .A3(new_n280_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n879_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n555_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n232_), .ZN(G1344gat));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n755_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n233_), .ZN(G1345gat));
  NOR2_X1   g720(.A1(new_n917_), .A2(new_n680_), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT61), .B(G155gat), .Z(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1346gat));
  NOR3_X1   g723(.A1(new_n917_), .A2(new_n225_), .A3(new_n666_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n916_), .A2(new_n681_), .A3(new_n879_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n225_), .B2(new_n926_), .ZN(G1347gat));
  INV_X1    g726(.A(new_n878_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n694_), .A2(new_n386_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n554_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT120), .ZN(new_n931_));
  OAI21_X1  g730(.A(G169gat), .B1(new_n928_), .B2(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT62), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n878_), .B2(new_n929_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n929_), .ZN(new_n936_));
  NOR4_X1   g735(.A1(new_n888_), .A2(KEYINPUT121), .A3(new_n281_), .A4(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n935_), .A2(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n554_), .B1(new_n407_), .B2(new_n404_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n933_), .B1(new_n938_), .B2(new_n939_), .ZN(G1348gat));
  OAI211_X1 g739(.A(new_n286_), .B(new_n623_), .C1(new_n935_), .C2(new_n937_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n878_), .A2(new_n623_), .A3(new_n929_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(G176gat), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n941_), .A2(KEYINPUT122), .A3(new_n943_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1349gat));
  INV_X1    g747(.A(new_n300_), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n637_), .B(new_n949_), .C1(new_n935_), .C2(new_n937_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n878_), .A2(new_n637_), .A3(new_n929_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(new_n409_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n950_), .A2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n950_), .A2(KEYINPUT123), .A3(new_n952_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n955_), .A2(new_n956_), .ZN(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n938_), .B2(new_n666_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n303_), .A2(new_n398_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n681_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n958_), .B1(new_n959_), .B2(new_n960_), .ZN(G1351gat));
  NAND2_X1  g760(.A1(new_n871_), .A2(new_n877_), .ZN(new_n962_));
  NAND4_X1  g761(.A1(new_n962_), .A2(new_n517_), .A3(new_n499_), .A4(new_n695_), .ZN(new_n963_));
  INV_X1    g762(.A(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(new_n554_), .ZN(new_n965_));
  OAI21_X1  g764(.A(KEYINPUT124), .B1(new_n965_), .B2(new_n206_), .ZN(new_n966_));
  OR4_X1    g765(.A1(KEYINPUT124), .A2(new_n963_), .A3(new_n206_), .A4(new_n555_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n965_), .A2(new_n206_), .ZN(new_n968_));
  AND3_X1   g767(.A1(new_n966_), .A2(new_n967_), .A3(new_n968_), .ZN(G1352gat));
  NAND2_X1  g768(.A1(new_n964_), .A2(new_n623_), .ZN(new_n970_));
  OAI22_X1  g769(.A1(new_n963_), .A2(new_n755_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n971_));
  NAND2_X1  g770(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n972_));
  MUX2_X1   g771(.A(new_n970_), .B(new_n971_), .S(new_n972_), .Z(G1353gat));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n974_), .A2(new_n630_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n976_));
  NAND4_X1  g775(.A1(new_n964_), .A2(new_n637_), .A3(new_n975_), .A4(new_n976_), .ZN(new_n977_));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n977_), .A2(new_n978_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n963_), .A2(new_n680_), .ZN(new_n980_));
  OR2_X1    g779(.A1(new_n980_), .A2(new_n975_), .ZN(new_n981_));
  NAND4_X1  g780(.A1(new_n980_), .A2(KEYINPUT126), .A3(new_n975_), .A4(new_n976_), .ZN(new_n982_));
  AND3_X1   g781(.A1(new_n979_), .A2(new_n981_), .A3(new_n982_), .ZN(G1354gat));
  NAND3_X1  g782(.A1(new_n964_), .A2(KEYINPUT127), .A3(new_n681_), .ZN(new_n984_));
  INV_X1    g783(.A(G218gat), .ZN(new_n985_));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986_));
  OAI21_X1  g785(.A(new_n986_), .B1(new_n963_), .B2(new_n661_), .ZN(new_n987_));
  NAND3_X1  g786(.A1(new_n984_), .A2(new_n985_), .A3(new_n987_), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n964_), .A2(G218gat), .A3(new_n665_), .ZN(new_n989_));
  AND2_X1   g788(.A1(new_n988_), .A2(new_n989_), .ZN(G1355gat));
endmodule


