//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n595_, new_n596_, new_n597_, new_n598_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_;
  NAND2_X1  g000(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT75), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n206_), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n205_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT66), .ZN(new_n213_));
  OR2_X1    g012(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n210_), .A2(new_n213_), .A3(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT65), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n221_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(G92gat), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n223_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT67), .B1(new_n218_), .B2(new_n228_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT66), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT66), .B1(new_n211_), .B2(new_n212_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(new_n224_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n220_), .A2(new_n222_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n232_), .A2(new_n235_), .A3(new_n236_), .A4(new_n217_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n229_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G85gat), .B(G92gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(KEYINPUT68), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  OR3_X1    g044(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n240_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n250_));
  NOR3_X1   g049(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n243_), .A2(new_n244_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n239_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT8), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n250_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n210_), .A2(new_n253_), .A3(new_n246_), .A4(new_n213_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(new_n255_), .A3(new_n240_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n249_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G29gat), .B(G36gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G43gat), .B(G50gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n238_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT73), .Z(new_n264_));
  NAND2_X1  g063(.A1(new_n238_), .A2(new_n259_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n262_), .B(KEYINPUT15), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT35), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G232gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT34), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n265_), .A2(new_n266_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n264_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n270_), .A2(new_n267_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n264_), .B(new_n271_), .C1(new_n267_), .C2(new_n270_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G190gat), .B(G218gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G134gat), .B(G162gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n279_), .B(KEYINPUT36), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n279_), .A2(KEYINPUT36), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n274_), .A2(new_n282_), .A3(new_n275_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n204_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n288_), .A3(new_n203_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G127gat), .B(G155gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT16), .ZN(new_n292_));
  XOR2_X1   g091(.A(G183gat), .B(G211gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT78), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT17), .Z(new_n296_));
  XNOR2_X1  g095(.A(G15gat), .B(G22gat), .ZN(new_n297_));
  INV_X1    g096(.A(G1gat), .ZN(new_n298_));
  INV_X1    g097(.A(G8gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT14), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G8gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G231gat), .A2(G233gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G57gat), .B(G64gat), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n306_), .A2(KEYINPUT11), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(KEYINPUT11), .ZN(new_n308_));
  XOR2_X1   g107(.A(G71gat), .B(G78gat), .Z(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n308_), .A2(new_n309_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n305_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT77), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n313_), .A2(KEYINPUT77), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n296_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n317_));
  OR3_X1    g116(.A1(new_n313_), .A2(new_n294_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n290_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT79), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n303_), .B(new_n262_), .Z(new_n323_));
  NAND2_X1  g122(.A1(G229gat), .A2(G233gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n266_), .A2(new_n303_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n303_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n327_), .B2(new_n262_), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n323_), .A2(new_n325_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G113gat), .B(G141gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(G169gat), .B(G197gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n329_), .B(new_n332_), .Z(new_n333_));
  INV_X1    g132(.A(KEYINPUT27), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT19), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n338_), .A2(KEYINPUT23), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G183gat), .ZN(new_n342_));
  INV_X1    g141(.A(G190gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT84), .B1(new_n341_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(G176gat), .B1(KEYINPUT83), .B2(KEYINPUT22), .ZN(new_n346_));
  INV_X1    g145(.A(G169gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n346_), .A2(new_n347_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n345_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n341_), .A2(KEYINPUT84), .A3(new_n344_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n340_), .A2(new_n337_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(KEYINPUT23), .B2(new_n337_), .ZN(new_n354_));
  MUX2_X1   g153(.A(new_n353_), .B(new_n354_), .S(KEYINPUT82), .Z(new_n355_));
  NOR2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT80), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT24), .ZN(new_n358_));
  INV_X1    g157(.A(G176gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n347_), .A2(new_n359_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT25), .B(G183gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT26), .B(G190gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n357_), .A2(new_n358_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n355_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G197gat), .B(G204gat), .Z(new_n367_));
  OR2_X1    g166(.A1(new_n367_), .A2(KEYINPUT21), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(KEYINPUT21), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n369_), .A2(new_n370_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n352_), .A2(new_n366_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n355_), .A2(new_n344_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G169gat), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n360_), .B1(new_n377_), .B2(new_n359_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n365_), .A2(new_n341_), .A3(KEYINPUT94), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n365_), .A2(new_n341_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT94), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n364_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n374_), .B1(new_n379_), .B2(new_n384_), .ZN(new_n385_));
  OAI211_X1 g184(.A(KEYINPUT20), .B(new_n375_), .C1(new_n385_), .C2(KEYINPUT95), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n385_), .A2(KEYINPUT95), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n336_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n352_), .A2(new_n366_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n373_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n379_), .A2(new_n374_), .A3(new_n384_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(KEYINPUT20), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n392_), .A2(new_n336_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT18), .ZN(new_n395_));
  XOR2_X1   g194(.A(G64gat), .B(G92gat), .Z(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n388_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n388_), .B2(new_n393_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n334_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n388_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n385_), .A2(KEYINPUT95), .ZN(new_n402_));
  INV_X1    g201(.A(new_n336_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n385_), .A2(KEYINPUT95), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n375_), .A2(KEYINPUT20), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n392_), .A2(new_n336_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(KEYINPUT27), .B(new_n401_), .C1(new_n408_), .C2(new_n397_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n400_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(G141gat), .ZN(new_n411_));
  INV_X1    g210(.A(G148gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n411_), .A2(new_n412_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G141gat), .A2(G148gat), .ZN(new_n418_));
  AOI22_X1  g217(.A1(KEYINPUT1), .A2(new_n417_), .B1(new_n418_), .B2(KEYINPUT87), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT1), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n413_), .A2(KEYINPUT3), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT89), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n414_), .A2(KEYINPUT2), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT3), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n431_), .B2(new_n418_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n427_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n423_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT90), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n424_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(KEYINPUT90), .A3(new_n423_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT28), .B1(new_n438_), .B2(KEYINPUT29), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT28), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n436_), .A2(new_n440_), .A3(new_n441_), .A4(new_n437_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G22gat), .B(G50gat), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n439_), .B2(new_n442_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT93), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n438_), .A2(KEYINPUT29), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(KEYINPUT92), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n441_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n373_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  OAI211_X1 g250(.A(G228gat), .B(G233gat), .C1(new_n448_), .C2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n447_), .A2(KEYINPUT91), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n374_), .B1(G228gat), .B2(G233gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G78gat), .B(G106gat), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n452_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n452_), .B2(new_n457_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n446_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n452_), .A2(new_n457_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n458_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n439_), .A2(new_n442_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n443_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT93), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n446_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n452_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n464_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n462_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n410_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G127gat), .B(G134gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G113gat), .B(G120gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n438_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n436_), .A2(new_n480_), .A3(new_n437_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(KEYINPUT4), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT96), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n482_), .B(new_n484_), .C1(KEYINPUT4), .C2(new_n479_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n479_), .A2(new_n481_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n483_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G1gat), .B(G29gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G57gat), .B(G85gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n490_), .B(new_n491_), .Z(new_n492_));
  NAND3_X1  g291(.A1(new_n485_), .A2(new_n487_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT98), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n485_), .A2(new_n487_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT98), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n485_), .A2(new_n487_), .A3(new_n498_), .A4(new_n492_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n494_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G71gat), .B(G99gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(G43gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G227gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(G15gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n502_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n389_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT85), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n509_), .B2(new_n508_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n509_), .A3(new_n506_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n478_), .B(KEYINPUT31), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(KEYINPUT86), .A3(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n513_), .A2(KEYINPUT86), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n514_), .B1(new_n513_), .B2(KEYINPUT86), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n475_), .A2(new_n500_), .A3(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n497_), .A2(new_n499_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n521_), .A2(new_n400_), .A3(new_n409_), .A4(new_n494_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(new_n474_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n462_), .A2(new_n473_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n398_), .A2(new_n399_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT33), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n493_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n493_), .A2(new_n526_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n492_), .B1(new_n486_), .B2(new_n484_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n482_), .B1(KEYINPUT4), .B2(new_n479_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n483_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n525_), .A2(new_n527_), .A3(new_n528_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n397_), .A2(KEYINPUT32), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n388_), .A2(new_n393_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n534_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n500_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n524_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n519_), .B1(new_n523_), .B2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n520_), .B1(new_n540_), .B2(KEYINPUT99), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT99), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n542_), .B(new_n519_), .C1(new_n523_), .C2(new_n539_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n333_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G230gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n238_), .A2(new_n259_), .A3(new_n312_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n312_), .B1(new_n238_), .B2(new_n259_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n546_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT70), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G120gat), .B(G148gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(G176gat), .B(G204gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(KEYINPUT71), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n547_), .A2(new_n545_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  INV_X1    g359(.A(new_n312_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n265_), .B2(new_n561_), .ZN(new_n562_));
  AOI211_X1 g361(.A(KEYINPUT12), .B(new_n312_), .C1(new_n238_), .C2(new_n259_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n559_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n552_), .A2(new_n558_), .A3(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n558_), .B1(new_n552_), .B2(new_n565_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT13), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n322_), .A2(new_n544_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n298_), .A3(new_n500_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT38), .ZN(new_n572_));
  INV_X1    g371(.A(new_n333_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(new_n319_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT100), .Z(new_n576_));
  XOR2_X1   g375(.A(new_n284_), .B(KEYINPUT101), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n500_), .ZN(new_n581_));
  OAI21_X1  g380(.A(G1gat), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT102), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n572_), .A2(new_n583_), .ZN(G1324gat));
  INV_X1    g383(.A(new_n410_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n570_), .A2(new_n299_), .A3(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G8gat), .B1(new_n580_), .B2(new_n410_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n587_), .A2(KEYINPUT39), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(KEYINPUT39), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n586_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT40), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT40), .B(new_n586_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(G1325gat));
  OAI21_X1  g393(.A(G15gat), .B1(new_n580_), .B2(new_n519_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT41), .Z(new_n596_));
  INV_X1    g395(.A(new_n519_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n570_), .A2(new_n504_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(G1326gat));
  OAI21_X1  g398(.A(G22gat), .B1(new_n580_), .B2(new_n474_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT42), .ZN(new_n601_));
  INV_X1    g400(.A(G22gat), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n570_), .A2(new_n602_), .A3(new_n524_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(G1327gat));
  NAND2_X1  g403(.A1(new_n285_), .A2(new_n319_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT103), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n569_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n544_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(G29gat), .B1(new_n611_), .B2(new_n500_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n574_), .A2(new_n320_), .ZN(new_n613_));
  AOI211_X1 g412(.A(KEYINPUT43), .B(new_n290_), .C1(new_n541_), .C2(new_n543_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n540_), .A2(KEYINPUT99), .ZN(new_n616_));
  INV_X1    g415(.A(new_n520_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n543_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n287_), .A2(new_n289_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n613_), .B1(new_n614_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT44), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(KEYINPUT44), .B(new_n613_), .C1(new_n614_), .C2(new_n620_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n500_), .A2(G29gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n612_), .B1(new_n625_), .B2(new_n626_), .ZN(G1328gat));
  INV_X1    g426(.A(KEYINPUT46), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(KEYINPUT104), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n623_), .A2(new_n585_), .A3(new_n624_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(G36gat), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n410_), .A2(G36gat), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n618_), .A2(new_n609_), .A3(new_n573_), .A4(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT45), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT45), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n544_), .A2(new_n636_), .A3(new_n609_), .A4(new_n633_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n635_), .A2(new_n637_), .B1(KEYINPUT104), .B2(new_n628_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n630_), .B1(new_n632_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  AOI211_X1 g439(.A(new_n629_), .B(new_n640_), .C1(new_n631_), .C2(G36gat), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n639_), .A2(new_n641_), .ZN(G1329gat));
  NAND4_X1  g441(.A1(new_n623_), .A2(G43gat), .A3(new_n597_), .A4(new_n624_), .ZN(new_n643_));
  INV_X1    g442(.A(G43gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n610_), .B2(new_n519_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g446(.A(G50gat), .B1(new_n611_), .B2(new_n524_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n524_), .A2(G50gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n625_), .B2(new_n649_), .ZN(G1331gat));
  AND2_X1   g449(.A1(new_n322_), .A2(new_n608_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n573_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G57gat), .B1(new_n655_), .B2(new_n500_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n319_), .A2(new_n573_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n579_), .A2(new_n608_), .A3(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n581_), .A2(KEYINPUT106), .ZN(new_n659_));
  MUX2_X1   g458(.A(KEYINPUT106), .B(new_n659_), .S(G57gat), .Z(new_n660_));
  AOI21_X1  g459(.A(new_n656_), .B1(new_n658_), .B2(new_n660_), .ZN(G1332gat));
  INV_X1    g460(.A(G64gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n658_), .B2(new_n585_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT48), .Z(new_n664_));
  INV_X1    g463(.A(new_n655_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n585_), .A2(new_n662_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT107), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n664_), .B1(new_n665_), .B2(new_n667_), .ZN(G1333gat));
  INV_X1    g467(.A(G71gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n655_), .A2(new_n669_), .A3(new_n597_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n658_), .B2(new_n597_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT49), .Z(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1334gat));
  INV_X1    g472(.A(G78gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n655_), .A2(new_n674_), .A3(new_n524_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n658_), .B2(new_n524_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT50), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1335gat));
  OR2_X1    g477(.A1(new_n614_), .A2(new_n620_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n569_), .A2(new_n573_), .A3(new_n320_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n225_), .A2(new_n226_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n681_), .A2(new_n581_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(G85gat), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n607_), .A2(new_n569_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n653_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n686_), .B2(new_n581_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n687_), .A2(new_n688_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n683_), .B1(new_n689_), .B2(new_n690_), .ZN(G1336gat));
  INV_X1    g490(.A(new_n686_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G92gat), .B1(new_n692_), .B2(new_n585_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT109), .ZN(new_n694_));
  INV_X1    g493(.A(new_n681_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n585_), .A2(G92gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(G1337gat));
  OAI21_X1  g496(.A(G99gat), .B1(new_n681_), .B2(new_n519_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n597_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n686_), .A2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT110), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT51), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT51), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n701_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1338gat));
  NAND3_X1  g505(.A1(new_n692_), .A2(new_n215_), .A3(new_n524_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n524_), .B(new_n680_), .C1(new_n614_), .C2(new_n620_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(G106gat), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G106gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT53), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT53), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n707_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1339gat));
  NOR3_X1   g515(.A1(new_n475_), .A2(new_n581_), .A3(new_n519_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT57), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n329_), .A2(new_n332_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n332_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n324_), .B1(new_n327_), .B2(new_n262_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n326_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n719_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT56), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n557_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n547_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n564_), .A2(KEYINPUT55), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n559_), .B(new_n731_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n732_));
  AOI221_X4 g531(.A(new_n728_), .B1(new_n546_), .B2(new_n729_), .C1(new_n730_), .C2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n732_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n729_), .A2(new_n546_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT112), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n727_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n735_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n728_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n734_), .A2(KEYINPUT112), .A3(new_n735_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n557_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n741_), .B2(KEYINPUT56), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n552_), .A2(new_n565_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n557_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n573_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n725_), .B1(new_n742_), .B2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n718_), .B1(new_n747_), .B2(new_n285_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n557_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n726_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n745_), .B1(new_n751_), .B2(new_n737_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT57), .B(new_n284_), .C1(new_n752_), .C2(new_n725_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n737_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT113), .B(new_n727_), .C1(new_n733_), .C2(new_n736_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n751_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n744_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(new_n724_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(KEYINPUT58), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n619_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT58), .B1(new_n757_), .B2(new_n759_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n748_), .B(new_n753_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n763_), .A2(new_n319_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n569_), .A2(new_n657_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n290_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(new_n290_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n717_), .B1(new_n764_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT114), .ZN(new_n771_));
  INV_X1    g570(.A(new_n769_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n763_), .A2(new_n319_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n717_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n771_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(G113gat), .B1(new_n777_), .B2(new_n573_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n763_), .A2(KEYINPUT116), .A3(new_n319_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT116), .B1(new_n763_), .B2(new_n319_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n772_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT115), .B(KEYINPUT59), .Z(new_n782_));
  NOR4_X1   g581(.A1(new_n475_), .A2(new_n519_), .A3(new_n581_), .A4(new_n782_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n781_), .A2(new_n783_), .B1(new_n770_), .B2(KEYINPUT59), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n573_), .A2(G113gat), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT117), .Z(new_n786_));
  AOI21_X1  g585(.A(new_n778_), .B1(new_n784_), .B2(new_n786_), .ZN(G1340gat));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n608_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n784_), .A2(KEYINPUT118), .A3(new_n608_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(G120gat), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(G120gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n569_), .B2(KEYINPUT60), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n777_), .B(new_n794_), .C1(KEYINPUT60), .C2(new_n793_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n795_), .ZN(G1341gat));
  AOI21_X1  g595(.A(G127gat), .B1(new_n777_), .B2(new_n320_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n320_), .A2(G127gat), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT119), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n784_), .B2(new_n799_), .ZN(G1342gat));
  NAND2_X1  g599(.A1(new_n784_), .A2(new_n619_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G134gat), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n577_), .A2(G134gat), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n771_), .A2(new_n776_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(KEYINPUT120), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  INV_X1    g606(.A(G134gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n784_), .B2(new_n619_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n807_), .B1(new_n809_), .B2(new_n804_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n810_), .ZN(G1343gat));
  NOR2_X1   g610(.A1(new_n597_), .A2(new_n474_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n585_), .A2(new_n581_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n774_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n573_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n608_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g617(.A(KEYINPUT61), .B(G155gat), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n814_), .A2(new_n821_), .A3(new_n320_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n814_), .B2(new_n320_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n820_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n824_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(new_n822_), .A3(new_n819_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1346gat));
  AND3_X1   g627(.A1(new_n814_), .A2(G162gat), .A3(new_n619_), .ZN(new_n829_));
  AOI21_X1  g628(.A(G162gat), .B1(new_n814_), .B2(new_n578_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n831_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n829_), .B1(new_n832_), .B2(new_n833_), .ZN(G1347gat));
  AND2_X1   g633(.A1(new_n781_), .A2(new_n474_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n519_), .A2(new_n410_), .A3(new_n500_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n836_), .A2(new_n377_), .A3(new_n573_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n573_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n840_), .A2(KEYINPUT123), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(KEYINPUT123), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n524_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n781_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n839_), .B1(new_n844_), .B2(G169gat), .ZN(new_n845_));
  AOI211_X1 g644(.A(KEYINPUT62), .B(new_n347_), .C1(new_n781_), .C2(new_n843_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n838_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT124), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n849_), .B(new_n838_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(G1348gat));
  NAND4_X1  g650(.A1(new_n781_), .A2(new_n474_), .A3(new_n608_), .A4(new_n836_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n359_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n524_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n854_), .A2(G176gat), .A3(new_n608_), .A4(new_n836_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT125), .ZN(G1349gat));
  NAND2_X1  g656(.A1(new_n835_), .A2(new_n836_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n858_), .A2(new_n362_), .A3(new_n319_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n854_), .A2(new_n320_), .A3(new_n836_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n342_), .B2(new_n860_), .ZN(G1350gat));
  OAI21_X1  g660(.A(G190gat), .B1(new_n858_), .B2(new_n290_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n578_), .A2(new_n363_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n858_), .B2(new_n863_), .ZN(G1351gat));
  NAND4_X1  g663(.A1(new_n774_), .A2(new_n581_), .A3(new_n585_), .A4(new_n812_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n333_), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g666(.A1(new_n865_), .A2(new_n569_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT126), .B(G204gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1353gat));
  AOI21_X1  g669(.A(new_n319_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT127), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n865_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1354gat));
  OAI21_X1  g674(.A(G218gat), .B1(new_n865_), .B2(new_n290_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n577_), .A2(G218gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n865_), .B2(new_n877_), .ZN(G1355gat));
endmodule


