//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202_));
  INV_X1    g001(.A(G134gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G127gat), .ZN(new_n204_));
  INV_X1    g003(.A(G127gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G134gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n202_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n204_), .A2(new_n206_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT84), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n202_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n210_), .A2(new_n215_), .A3(KEYINPUT85), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(KEYINPUT85), .B2(new_n210_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT31), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n227_), .ZN(new_n228_));
  OR3_X1    g027(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n223_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(KEYINPUT81), .A2(KEYINPUT26), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT81), .A2(KEYINPUT26), .ZN(new_n232_));
  OAI21_X1  g031(.A(G190gat), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G183gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT79), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G183gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT78), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT78), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G183gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n243_), .A3(KEYINPUT25), .ZN(new_n244_));
  OR2_X1    g043(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT26), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n244_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n230_), .B1(new_n239_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n227_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n224_), .A2(KEYINPUT22), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT22), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G169gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT82), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(G176gat), .B1(new_n252_), .B2(KEYINPUT82), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n251_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n245_), .A2(new_n241_), .A3(new_n243_), .A4(new_n246_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n220_), .A2(new_n222_), .A3(KEYINPUT83), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n219_), .A2(new_n262_), .A3(KEYINPUT23), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n250_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G71gat), .B(G99gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G43gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n266_), .B(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G227gat), .A2(G233gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n270_), .B(G15gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT30), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n269_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT86), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n218_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(KEYINPUT86), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n273_), .A2(KEYINPUT86), .A3(new_n218_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT88), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(KEYINPUT88), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290_));
  INV_X1    g089(.A(G141gat), .ZN(new_n291_));
  INV_X1    g090(.A(G148gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT2), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT89), .B1(new_n289_), .B2(new_n298_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n287_), .A2(new_n288_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n284_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n294_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n283_), .B1(new_n281_), .B2(KEYINPUT1), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT87), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n283_), .A2(KEYINPUT1), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n307_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n217_), .B1(new_n304_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n284_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n289_), .A2(KEYINPUT89), .A3(new_n298_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n301_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n210_), .A2(new_n215_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n313_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n314_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n314_), .A2(KEYINPUT4), .A3(new_n321_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n320_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT4), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n217_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n322_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n323_), .B1(new_n324_), .B2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G1gat), .B(G29gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G85gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT0), .B(G57gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n334_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n323_), .B(new_n336_), .C1(new_n324_), .C2(new_n329_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G8gat), .B(G36gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT18), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n257_), .A2(new_n258_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n343_), .A2(new_n264_), .A3(new_n227_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n223_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n233_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n346_));
  XOR2_X1   g145(.A(KEYINPUT80), .B(G190gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT78), .B(G183gat), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n347_), .A2(KEYINPUT26), .B1(new_n348_), .B2(KEYINPUT25), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n351_));
  INV_X1    g150(.A(G211gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n352_), .B2(G218gat), .ZN(new_n353_));
  INV_X1    g152(.A(G218gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(G211gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G197gat), .ZN(new_n357_));
  INV_X1    g156(.A(G204gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G197gat), .A2(G204gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(KEYINPUT21), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT21), .ZN(new_n362_));
  AND2_X1   g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n356_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n363_), .A2(new_n364_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n367_), .B(KEYINPUT21), .C1(new_n355_), .C2(new_n353_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n366_), .A2(KEYINPUT91), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT91), .B1(new_n366_), .B2(new_n368_), .ZN(new_n370_));
  OAI22_X1  g169(.A1(new_n344_), .A2(new_n350_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT96), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT22), .B(G169gat), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n251_), .B1(new_n373_), .B2(new_n225_), .ZN(new_n374_));
  INV_X1    g173(.A(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n240_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n223_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n240_), .A2(KEYINPUT25), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n235_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n248_), .A2(G190gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n375_), .A2(KEYINPUT26), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT95), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n375_), .A2(KEYINPUT26), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n248_), .A2(G190gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT95), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n380_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n261_), .A2(new_n228_), .A3(new_n263_), .A4(new_n229_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n378_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n366_), .A2(new_n368_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n372_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n380_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n386_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n261_), .A2(new_n263_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n228_), .A2(new_n229_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n366_), .A2(new_n368_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT96), .A4(new_n378_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n371_), .A2(new_n392_), .A3(KEYINPUT20), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT19), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT91), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n391_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n366_), .A2(new_n368_), .A3(KEYINPUT91), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n250_), .A4(new_n265_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n390_), .A2(new_n391_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n410_), .A2(KEYINPUT20), .A3(new_n404_), .A4(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT98), .B1(new_n406_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n399_), .A2(new_n400_), .A3(new_n378_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n369_), .A2(new_n370_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n346_), .A2(new_n349_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n416_), .A2(new_n230_), .B1(new_n259_), .B2(new_n264_), .ZN(new_n417_));
  OAI211_X1 g216(.A(KEYINPUT20), .B(new_n414_), .C1(new_n415_), .C2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n404_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n410_), .A2(KEYINPUT20), .A3(new_n405_), .A4(new_n411_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT32), .B(new_n342_), .C1(new_n413_), .C2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n406_), .A2(new_n412_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n342_), .A2(KEYINPUT32), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(KEYINPUT98), .A3(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n338_), .A2(new_n422_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n342_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n406_), .A2(new_n412_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n406_), .B2(new_n412_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n314_), .A2(new_n321_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n334_), .B1(new_n431_), .B2(new_n322_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT97), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI211_X1 g233(.A(KEYINPUT97), .B(new_n334_), .C1(new_n431_), .C2(new_n322_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n322_), .B(new_n327_), .C1(new_n431_), .C2(new_n326_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n337_), .A2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n328_), .B(new_n327_), .C1(new_n431_), .C2(new_n326_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n440_), .A2(KEYINPUT33), .A3(new_n323_), .A4(new_n336_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n430_), .A2(new_n437_), .A3(new_n439_), .A4(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n426_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT94), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT28), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n304_), .A2(new_n313_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT29), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NOR4_X1   g249(.A1(new_n304_), .A2(KEYINPUT28), .A3(new_n313_), .A4(KEYINPUT29), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G22gat), .B(G50gat), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT28), .B1(new_n325_), .B2(KEYINPUT29), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n448_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n446_), .B1(new_n453_), .B2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n449_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n408_), .A2(new_n409_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G228gat), .A2(G233gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT92), .B1(new_n459_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT29), .B1(new_n304_), .B2(new_n313_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT92), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n461_), .A4(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n461_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n459_), .B2(new_n400_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(KEYINPUT93), .B(new_n468_), .C1(new_n459_), .C2(new_n400_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n467_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n452_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n455_), .A2(new_n456_), .A3(new_n454_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n444_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n458_), .A2(new_n473_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n473_), .B1(new_n458_), .B2(new_n477_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n443_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n479_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n458_), .A2(new_n473_), .A3(new_n477_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n338_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n423_), .A2(new_n342_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n406_), .A2(new_n412_), .A3(new_n427_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT27), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n342_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT27), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n429_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n484_), .A2(new_n485_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n280_), .B1(new_n481_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n490_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT99), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n497_), .B1(new_n460_), .B2(new_n266_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n405_), .B1(new_n498_), .B2(new_n414_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n420_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n427_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n412_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(new_n405_), .B2(new_n402_), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT27), .B(new_n501_), .C1(new_n503_), .C2(new_n427_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n495_), .A2(new_n496_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n496_), .B1(new_n495_), .B2(new_n504_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n480_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT100), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT99), .B1(new_n488_), .B2(new_n491_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n495_), .A2(new_n496_), .A3(new_n504_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT100), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n480_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n278_), .A2(new_n279_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(new_n338_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n494_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G15gat), .B(G22gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT70), .B(G1gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(G8gat), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n520_), .B2(KEYINPUT14), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT71), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G8gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n521_), .A2(KEYINPUT71), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n521_), .A2(KEYINPUT71), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n523_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G29gat), .B(G36gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT68), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G43gat), .B(G50gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n525_), .A2(new_n528_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(KEYINPUT75), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n538_), .A2(new_n540_), .A3(G229gat), .A4(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n532_), .B(KEYINPUT15), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n525_), .A2(new_n528_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT76), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n537_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G169gat), .B(G197gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n548_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT77), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n541_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n548_), .A2(KEYINPUT77), .A3(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n517_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G85gat), .B(G92gat), .Z(new_n560_));
  NOR2_X1   g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT6), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n560_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT65), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT8), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT10), .B(G99gat), .Z(new_n572_));
  INV_X1    g371(.A(G106gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT64), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(G85gat), .ZN(new_n577_));
  INV_X1    g376(.A(G92gat), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT9), .ZN(new_n579_));
  AOI211_X1 g378(.A(new_n579_), .B(new_n566_), .C1(KEYINPUT9), .C2(new_n560_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n571_), .A2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n567_), .A2(new_n568_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n569_), .A2(new_n583_), .A3(new_n570_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT66), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  OR3_X1    g384(.A1(new_n569_), .A2(new_n583_), .A3(new_n570_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT66), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n570_), .A2(new_n569_), .B1(new_n576_), .B2(new_n580_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G57gat), .B(G64gat), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT11), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(KEYINPUT11), .ZN(new_n592_));
  XOR2_X1   g391(.A(G71gat), .B(G78gat), .Z(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT12), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n585_), .A2(new_n589_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n586_), .A2(new_n596_), .A3(new_n588_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n597_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .A4(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n602_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(G230gat), .A3(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT5), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n610_), .B(new_n611_), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n606_), .A2(new_n608_), .A3(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT67), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n606_), .A2(new_n608_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n612_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT13), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n615_), .A2(KEYINPUT13), .A3(new_n617_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(KEYINPUT69), .A2(KEYINPUT37), .ZN(new_n623_));
  NAND2_X1  g422(.A1(KEYINPUT69), .A2(KEYINPUT37), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT36), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n585_), .A2(new_n589_), .A3(new_n542_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT34), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(KEYINPUT35), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n582_), .A2(new_n584_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n633_), .B2(new_n532_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(KEYINPUT35), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n629_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n635_), .B1(new_n629_), .B2(new_n634_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n628_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n638_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n627_), .A2(KEYINPUT36), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n636_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n623_), .B(new_n624_), .C1(new_n640_), .C2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n642_), .A3(new_n636_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n639_), .A2(new_n645_), .A3(KEYINPUT69), .A4(KEYINPUT37), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G127gat), .B(G155gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT16), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G183gat), .B(G211gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(KEYINPUT73), .B(KEYINPUT17), .Z(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT74), .Z(new_n654_));
  NAND2_X1  g453(.A1(G231gat), .A2(G233gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n596_), .B(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n543_), .B(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT72), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n659_), .B1(new_n658_), .B2(new_n657_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n651_), .B(KEYINPUT17), .Z(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n647_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n559_), .A2(new_n622_), .A3(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n665_), .A2(new_n485_), .A3(new_n519_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n666_), .A2(KEYINPUT38), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(KEYINPUT38), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n640_), .A2(new_n643_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n517_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n558_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n663_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n622_), .A4(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G1gat), .B1(new_n673_), .B2(new_n485_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n667_), .A2(new_n668_), .A3(new_n674_), .ZN(G1324gat));
  OAI21_X1  g474(.A(G8gat), .B1(new_n673_), .B2(new_n511_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(KEYINPUT39), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n665_), .A2(G8gat), .A3(new_n511_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n676_), .A2(new_n677_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(KEYINPUT39), .A3(new_n678_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1325gat));
  OAI21_X1  g485(.A(G15gat), .B1(new_n673_), .B2(new_n515_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT41), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n665_), .A2(G15gat), .A3(new_n515_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1326gat));
  OAI21_X1  g489(.A(G22gat), .B1(new_n673_), .B2(new_n480_), .ZN(new_n691_));
  XOR2_X1   g490(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n480_), .A2(G22gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n665_), .B2(new_n694_), .ZN(G1327gat));
  AND2_X1   g494(.A1(new_n644_), .A2(new_n646_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n517_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n280_), .A2(new_n485_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n508_), .B2(new_n513_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n698_), .B(new_n647_), .C1(new_n700_), .C2(new_n494_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n620_), .A2(new_n671_), .A3(new_n621_), .A4(new_n663_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT44), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n706_), .B(new_n703_), .C1(new_n697_), .C2(new_n701_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n338_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G29gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n708_), .B2(new_n338_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n511_), .A2(new_n512_), .A3(new_n480_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n512_), .B1(new_n511_), .B2(new_n480_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n516_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n494_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n669_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(new_n672_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n717_), .A2(new_n671_), .A3(new_n622_), .A4(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n485_), .A2(G29gat), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT104), .Z(new_n722_));
  OAI22_X1  g521(.A1(new_n711_), .A2(new_n712_), .B1(new_n720_), .B2(new_n722_), .ZN(G1328gat));
  AOI21_X1  g522(.A(new_n698_), .B1(new_n717_), .B2(new_n647_), .ZN(new_n724_));
  AOI211_X1 g523(.A(KEYINPUT43), .B(new_n696_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n704_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n706_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n511_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n702_), .A2(KEYINPUT44), .A3(new_n704_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n511_), .B(KEYINPUT106), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(G36gat), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n720_), .A2(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT45), .Z(new_n737_));
  NAND2_X1  g536(.A1(new_n731_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT105), .B1(new_n730_), .B2(G36gat), .ZN(new_n739_));
  OAI211_X1 g538(.A(KEYINPUT107), .B(KEYINPUT46), .C1(new_n738_), .C2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n705_), .A2(new_n707_), .A3(new_n511_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(new_n734_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(new_n731_), .A3(new_n737_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT46), .B1(new_n745_), .B2(KEYINPUT107), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n741_), .A2(new_n746_), .ZN(G1329gat));
  NOR3_X1   g546(.A1(new_n720_), .A2(G43gat), .A3(new_n515_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n708_), .A2(new_n280_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(G43gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g550(.A1(new_n720_), .A2(new_n480_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(G50gat), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n484_), .A2(G50gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n708_), .B2(new_n754_), .ZN(G1331gat));
  INV_X1    g554(.A(new_n622_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n664_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT108), .Z(new_n758_));
  NOR3_X1   g557(.A1(new_n758_), .A2(new_n517_), .A3(new_n671_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT109), .ZN(new_n760_));
  INV_X1    g559(.A(G57gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n338_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n622_), .A2(new_n671_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n670_), .A2(new_n672_), .A3(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G57gat), .B1(new_n764_), .B2(new_n485_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1332gat));
  INV_X1    g565(.A(G64gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n760_), .A2(new_n767_), .A3(new_n733_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G64gat), .B1(new_n764_), .B2(new_n732_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT48), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1333gat));
  NOR2_X1   g570(.A1(new_n515_), .A2(G71gat), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT110), .Z(new_n773_));
  NAND2_X1  g572(.A1(new_n760_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G71gat), .B1(new_n764_), .B2(new_n515_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT49), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1334gat));
  INV_X1    g576(.A(G78gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n760_), .A2(new_n778_), .A3(new_n484_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G78gat), .B1(new_n764_), .B2(new_n480_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT111), .Z(new_n781_));
  OR2_X1    g580(.A1(new_n781_), .A2(KEYINPUT50), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(KEYINPUT50), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n779_), .A2(new_n782_), .A3(new_n783_), .ZN(G1335gat));
  NAND4_X1  g583(.A1(new_n756_), .A2(new_n717_), .A3(new_n558_), .A4(new_n719_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n577_), .A3(new_n338_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n702_), .A2(new_n663_), .A3(new_n763_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(new_n338_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n787_), .B1(new_n789_), .B2(new_n577_), .ZN(G1336gat));
  NOR3_X1   g589(.A1(new_n785_), .A2(G92gat), .A3(new_n511_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n788_), .A2(new_n733_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G92gat), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT112), .ZN(G1337gat));
  INV_X1    g593(.A(G99gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n788_), .B2(new_n280_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n786_), .A2(new_n280_), .A3(new_n572_), .ZN(new_n797_));
  OAI22_X1  g596(.A1(new_n796_), .A2(new_n797_), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n798_));
  NAND2_X1  g597(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(G1338gat));
  NAND3_X1  g599(.A1(new_n786_), .A2(new_n573_), .A3(new_n484_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n788_), .A2(new_n484_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(G106gat), .ZN(new_n804_));
  AOI211_X1 g603(.A(KEYINPUT52), .B(new_n573_), .C1(new_n788_), .C2(new_n484_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(KEYINPUT114), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n622_), .A2(new_n558_), .A3(new_n664_), .A4(new_n809_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n622_), .A2(new_n558_), .A3(new_n664_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n538_), .A2(new_n540_), .A3(new_n546_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n536_), .A2(new_n546_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n551_), .B1(new_n815_), .B2(new_n544_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n615_), .A2(new_n555_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n606_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT115), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n606_), .A2(new_n819_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n600_), .A2(new_n602_), .A3(new_n605_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(G230gat), .A3(G233gat), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n606_), .A2(new_n825_), .A3(new_n819_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n821_), .A2(new_n822_), .A3(new_n824_), .A4(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(KEYINPUT56), .A3(new_n612_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n827_), .B2(new_n612_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(KEYINPUT116), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n612_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n831_), .A2(KEYINPUT116), .A3(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n818_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT58), .B(new_n818_), .C1(new_n830_), .C2(new_n833_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n647_), .A3(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n556_), .A2(new_n615_), .A3(new_n557_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n831_), .A2(new_n832_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n828_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n618_), .A2(new_n555_), .A3(new_n817_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n718_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT57), .B(new_n718_), .C1(new_n841_), .C2(new_n843_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n838_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n813_), .B1(new_n848_), .B2(new_n663_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n514_), .A2(new_n338_), .A3(new_n280_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(G113gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n671_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n850_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n846_), .A2(new_n847_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n672_), .B1(new_n857_), .B2(new_n838_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT59), .B(new_n856_), .C1(new_n858_), .C2(new_n813_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n558_), .B1(new_n855_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n853_), .B1(new_n860_), .B2(new_n852_), .ZN(G1340gat));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n622_), .B2(KEYINPUT60), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n851_), .B(new_n863_), .C1(KEYINPUT60), .C2(new_n862_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n622_), .B1(new_n855_), .B2(new_n859_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866_));
  OAI21_X1  g665(.A(G120gat), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  AOI211_X1 g666(.A(KEYINPUT118), .B(new_n622_), .C1(new_n855_), .C2(new_n859_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n867_), .B2(new_n868_), .ZN(G1341gat));
  AOI21_X1  g668(.A(G127gat), .B1(new_n851_), .B2(new_n672_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n855_), .A2(new_n859_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n663_), .A2(KEYINPUT119), .ZN(new_n872_));
  MUX2_X1   g671(.A(KEYINPUT119), .B(new_n872_), .S(G127gat), .Z(new_n873_));
  AOI21_X1  g672(.A(new_n870_), .B1(new_n871_), .B2(new_n873_), .ZN(G1342gat));
  NAND3_X1  g673(.A1(new_n851_), .A2(new_n203_), .A3(new_n669_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n696_), .B1(new_n855_), .B2(new_n859_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n203_), .ZN(G1343gat));
  NOR3_X1   g676(.A1(new_n733_), .A2(new_n485_), .A3(new_n480_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n515_), .B(new_n878_), .C1(new_n858_), .C2(new_n813_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n558_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n291_), .ZN(G1344gat));
  OAI21_X1  g680(.A(KEYINPUT121), .B1(new_n879_), .B2(new_n622_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n849_), .A2(new_n280_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n883_), .A2(new_n884_), .A3(new_n756_), .A4(new_n878_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT120), .B(G148gat), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n882_), .A2(new_n885_), .A3(new_n887_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1345gat));
  NOR2_X1   g690(.A1(new_n879_), .A2(new_n663_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT61), .B(G155gat), .Z(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  INV_X1    g693(.A(G162gat), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n879_), .A2(new_n895_), .A3(new_n696_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n879_), .B2(new_n718_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  OAI211_X1 g698(.A(KEYINPUT122), .B(new_n895_), .C1(new_n879_), .C2(new_n718_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n896_), .B1(new_n899_), .B2(new_n900_), .ZN(G1347gat));
  INV_X1    g700(.A(new_n849_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n732_), .A2(new_n699_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n671_), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT123), .Z(new_n905_));
  NAND3_X1  g704(.A1(new_n902_), .A2(new_n480_), .A3(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n906_), .A2(new_n907_), .A3(G169gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n906_), .B2(G169gat), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n480_), .B(new_n903_), .C1(new_n858_), .C2(new_n813_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n671_), .A2(new_n373_), .ZN(new_n911_));
  OAI22_X1  g710(.A1(new_n908_), .A2(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(G1348gat));
  NOR2_X1   g711(.A1(new_n910_), .A2(new_n622_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(new_n225_), .ZN(G1349gat));
  OR2_X1    g713(.A1(new_n910_), .A2(new_n663_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n393_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n348_), .B2(new_n915_), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n910_), .B2(new_n696_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n718_), .B1(new_n387_), .B2(new_n383_), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n902_), .A2(new_n480_), .A3(new_n903_), .A4(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT124), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n918_), .A2(new_n920_), .A3(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1351gat));
  NOR3_X1   g724(.A1(new_n732_), .A2(new_n338_), .A3(new_n480_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n883_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n558_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(new_n357_), .ZN(G1352gat));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n622_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(new_n358_), .ZN(G1353gat));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n663_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT125), .ZN(new_n934_));
  OAI221_X1 g733(.A(new_n932_), .B1(KEYINPUT63), .B2(G211gat), .C1(new_n927_), .C2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n927_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n932_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n932_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n934_), .A2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n936_), .A2(new_n937_), .A3(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n935_), .A2(new_n940_), .ZN(G1354gat));
  XNOR2_X1  g740(.A(KEYINPUT127), .B(G218gat), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n927_), .A2(new_n696_), .A3(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n936_), .A2(new_n669_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n944_), .B2(new_n942_), .ZN(G1355gat));
endmodule


