//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n207_), .B(KEYINPUT90), .Z(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G127gat), .B(G134gat), .ZN(new_n210_));
  INV_X1    g009(.A(G113gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G120gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n210_), .B(G113gat), .ZN(new_n214_));
  INV_X1    g013(.A(G120gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n220_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  OR2_X1    g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(KEYINPUT1), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n228_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n231_), .B1(new_n230_), .B2(new_n228_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n227_), .A2(KEYINPUT1), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n221_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(new_n218_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n229_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT91), .B(KEYINPUT4), .Z(new_n240_));
  NAND3_X1  g039(.A1(new_n217_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  OAI211_X1 g043(.A(KEYINPUT89), .B(new_n229_), .C1(new_n235_), .C2(new_n238_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n217_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n213_), .A2(new_n216_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(new_n243_), .A3(new_n239_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  AOI211_X1 g048(.A(new_n209_), .B(new_n242_), .C1(new_n249_), .C2(KEYINPUT4), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n208_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n206_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(KEYINPUT4), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(new_n208_), .A3(new_n241_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n251_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n206_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n252_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G71gat), .B(G99gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G15gat), .B(G43gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT24), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  MUX2_X1   g063(.A(new_n263_), .B(KEYINPUT24), .S(new_n264_), .Z(new_n265_));
  INV_X1    g064(.A(G183gat), .ZN(new_n266_));
  INV_X1    g065(.A(G190gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT23), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(new_n268_), .ZN(new_n272_));
  AND2_X1   g071(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n273_));
  NOR2_X1   g072(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT26), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT76), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT76), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT26), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n279_), .A3(G190gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT74), .B1(new_n281_), .B2(G183gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n275_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT25), .B(G183gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n284_), .A2(KEYINPUT74), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n265_), .B(new_n272_), .C1(new_n283_), .C2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n287_));
  INV_X1    g086(.A(G176gat), .ZN(new_n288_));
  AND2_X1   g087(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n269_), .B1(G183gat), .B2(G190gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(new_n271_), .B2(new_n268_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n273_), .A2(new_n274_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(G183gat), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n262_), .B(new_n291_), .C1(new_n293_), .C2(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n286_), .A2(new_n287_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n287_), .B1(new_n286_), .B2(new_n296_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n261_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n286_), .A2(new_n296_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT30), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n286_), .A2(new_n287_), .A3(new_n296_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n261_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G227gat), .A2(G233gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n305_), .B(KEYINPUT78), .Z(new_n306_));
  AND3_X1   g105(.A1(new_n299_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n299_), .B2(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT79), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n247_), .A2(KEYINPUT31), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n217_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n309_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n307_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n313_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n306_), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n297_), .A2(new_n298_), .A3(new_n261_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n303_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n299_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n315_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n260_), .B1(new_n314_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n313_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n259_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n239_), .A2(KEYINPUT29), .ZN(new_n327_));
  XOR2_X1   g126(.A(G22gat), .B(G50gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT28), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n327_), .B(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G78gat), .B(G106gat), .Z(new_n331_));
  INV_X1    g130(.A(G228gat), .ZN(new_n332_));
  INV_X1    g131(.A(G233gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n239_), .A2(KEYINPUT29), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G211gat), .A2(G218gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT21), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G211gat), .A2(G218gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(G211gat), .A2(G218gat), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n344_), .A2(new_n339_), .A3(KEYINPUT81), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n338_), .B(new_n343_), .C1(new_n345_), .C2(new_n341_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n342_), .ZN(new_n347_));
  OAI211_X1 g146(.A(KEYINPUT21), .B(new_n337_), .C1(new_n347_), .C2(KEYINPUT81), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n335_), .B1(new_n336_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT82), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n346_), .A2(KEYINPUT82), .A3(new_n348_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(new_n336_), .A3(new_n335_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n331_), .B1(new_n351_), .B2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n330_), .B1(new_n357_), .B2(KEYINPUT83), .ZN(new_n358_));
  INV_X1    g157(.A(new_n331_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n356_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n359_), .B1(new_n360_), .B2(new_n350_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n351_), .A2(new_n356_), .A3(new_n331_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n362_), .A3(new_n330_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT84), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n361_), .A2(new_n362_), .A3(KEYINPUT84), .A4(new_n330_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n258_), .B1(new_n326_), .B2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n368_), .A2(new_n369_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n372_), .A2(new_n365_), .A3(new_n325_), .A4(new_n322_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n346_), .A2(KEYINPUT82), .A3(new_n348_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT82), .B1(new_n346_), .B2(new_n348_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n300_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT85), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT19), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n272_), .B1(G183gat), .B2(G190gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT87), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n289_), .A2(new_n290_), .A3(KEYINPUT86), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT86), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT22), .ZN(new_n385_));
  INV_X1    g184(.A(G169gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n384_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n288_), .B1(new_n383_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n382_), .B1(new_n390_), .B2(new_n262_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT86), .B1(new_n289_), .B2(new_n290_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n387_), .A2(new_n384_), .A3(new_n388_), .ZN(new_n393_));
  AOI21_X1  g192(.A(G176gat), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n262_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n394_), .A2(KEYINPUT87), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n381_), .B1(new_n391_), .B2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(KEYINPUT26), .B(G190gat), .Z(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n293_), .B1(new_n284_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n265_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n349_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n353_), .A2(new_n354_), .A3(new_n296_), .A4(new_n286_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT85), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(KEYINPUT20), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n378_), .A2(new_n380_), .A3(new_n403_), .A4(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n349_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n397_), .A2(new_n408_), .A3(new_n401_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n355_), .A2(new_n300_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(KEYINPUT20), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n380_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT18), .B(G64gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G92gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n407_), .A2(new_n413_), .A3(new_n418_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT27), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(KEYINPUT88), .A3(new_n419_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT94), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n411_), .B2(new_n380_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n378_), .A2(new_n412_), .A3(new_n403_), .A4(new_n406_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n404_), .A2(KEYINPUT20), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n431_), .A2(KEYINPUT85), .B1(new_n402_), .B2(new_n349_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n432_), .A2(new_n427_), .A3(new_n412_), .A4(new_n406_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n418_), .A3(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(KEYINPUT27), .A3(new_n420_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n371_), .A2(new_n373_), .A3(new_n426_), .A4(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n419_), .A2(KEYINPUT32), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n430_), .A2(new_n438_), .A3(new_n433_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT95), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT95), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n430_), .A2(new_n441_), .A3(new_n438_), .A4(new_n433_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n414_), .A2(new_n437_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n414_), .A2(KEYINPUT93), .A3(new_n437_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n446_), .A2(new_n447_), .B1(new_n252_), .B2(new_n257_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n423_), .A2(new_n425_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n242_), .B1(new_n249_), .B2(KEYINPUT4), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n209_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n249_), .A2(new_n208_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n451_), .A2(new_n206_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n257_), .A2(KEYINPUT33), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n251_), .B1(new_n450_), .B2(new_n208_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n256_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n453_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n443_), .A2(new_n448_), .B1(new_n449_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n436_), .B1(new_n459_), .B2(new_n373_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462_));
  INV_X1    g261(.A(G1gat), .ZN(new_n463_));
  INV_X1    g262(.A(G8gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT14), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G1gat), .B(G8gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n466_), .B(new_n467_), .Z(new_n468_));
  XNOR2_X1  g267(.A(G57gat), .B(G64gat), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n469_), .A2(KEYINPUT11), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(KEYINPUT11), .ZN(new_n471_));
  XOR2_X1   g270(.A(G71gat), .B(G78gat), .Z(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n471_), .A2(new_n472_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n468_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G231gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT17), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT16), .B(G183gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(G211gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(G127gat), .B(G155gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  OR3_X1    g283(.A1(new_n479_), .A2(new_n480_), .A3(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(KEYINPUT17), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G50gat), .ZN(new_n489_));
  OR2_X1    g288(.A1(G29gat), .A2(G36gat), .ZN(new_n490_));
  INV_X1    g289(.A(G43gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G29gat), .A2(G36gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n491_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n489_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n490_), .A2(new_n492_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G43gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G50gat), .A3(new_n493_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n496_), .A2(KEYINPUT15), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT15), .B1(new_n496_), .B2(new_n499_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT8), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT7), .ZN(new_n505_));
  INV_X1    g304(.A(G99gat), .ZN(new_n506_));
  INV_X1    g305(.A(G106gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n508_), .A2(new_n511_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G85gat), .B(G92gat), .Z(new_n515_));
  AOI21_X1  g314(.A(new_n504_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n514_), .A2(new_n504_), .A3(new_n515_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT65), .B1(G85gat), .B2(G92gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n524_), .A2(G85gat), .A3(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n520_), .B(new_n523_), .C1(new_n526_), .C2(KEYINPUT9), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT10), .B(G99gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(G106gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n511_), .A2(new_n512_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n527_), .A2(new_n531_), .A3(KEYINPUT66), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT66), .B1(new_n527_), .B2(new_n531_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n519_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n494_), .A2(new_n489_), .A3(new_n495_), .ZN(new_n535_));
  AOI21_X1  g334(.A(G50gat), .B1(new_n498_), .B2(new_n493_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n517_), .A2(new_n518_), .B1(new_n527_), .B2(new_n531_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n503_), .A2(new_n534_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT34), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n539_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n542_), .A2(new_n543_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n539_), .A2(KEYINPUT35), .A3(new_n541_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(G134gat), .ZN(new_n552_));
  INV_X1    g351(.A(G162gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT36), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n554_), .B(KEYINPUT36), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n550_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n461_), .A2(new_n488_), .A3(new_n562_), .ZN(new_n563_));
  OR3_X1    g362(.A1(new_n502_), .A2(KEYINPUT72), .A3(new_n468_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n537_), .A2(KEYINPUT71), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n537_), .A2(KEYINPUT71), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n468_), .A3(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT72), .B1(new_n502_), .B2(new_n468_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n564_), .A2(new_n565_), .A3(new_n568_), .A4(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n565_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n568_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n468_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G169gat), .B(G197gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(G141gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT73), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n211_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n579_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n570_), .A2(new_n574_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n538_), .B(new_n475_), .Z(new_n585_));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT67), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n527_), .A2(new_n531_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n475_), .B1(new_n519_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n588_), .B1(new_n590_), .B2(KEYINPUT12), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT12), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT67), .B(new_n592_), .C1(new_n538_), .C2(new_n475_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n475_), .A2(new_n592_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n534_), .A2(new_n595_), .B1(new_n538_), .B2(new_n475_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n594_), .A2(KEYINPUT68), .A3(new_n586_), .A4(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n596_), .A2(new_n591_), .A3(new_n593_), .A4(new_n586_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT68), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n587_), .B1(new_n597_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT69), .B(G204gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT5), .B(G176gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n604_), .B(new_n605_), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT70), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n601_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT13), .ZN(new_n610_));
  INV_X1    g409(.A(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n601_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n609_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n601_), .A2(new_n608_), .ZN(new_n614_));
  AOI211_X1 g413(.A(new_n606_), .B(new_n587_), .C1(new_n597_), .C2(new_n600_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT13), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n584_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n563_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n258_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G1gat), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT97), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n558_), .A2(KEYINPUT37), .A3(new_n560_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n550_), .A2(new_n559_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n624_), .B2(new_n557_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n622_), .A2(new_n625_), .A3(new_n488_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n460_), .A2(new_n617_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(KEYINPUT38), .ZN(new_n629_));
  NOR4_X1   g428(.A1(new_n627_), .A2(G1gat), .A3(new_n619_), .A4(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(KEYINPUT38), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n621_), .A2(new_n632_), .ZN(G1324gat));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n634_));
  INV_X1    g433(.A(new_n618_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n426_), .A2(new_n435_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n637_), .B2(G8gat), .ZN(new_n638_));
  AOI211_X1 g437(.A(KEYINPUT39), .B(new_n464_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n464_), .ZN(new_n640_));
  OAI22_X1  g439(.A1(new_n638_), .A2(new_n639_), .B1(new_n627_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(G1325gat));
  INV_X1    g442(.A(new_n326_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G15gat), .B1(new_n618_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT41), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n627_), .A2(G15gat), .A3(new_n644_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1326gat));
  INV_X1    g447(.A(new_n370_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G22gat), .B1(new_n618_), .B2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT42), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n649_), .A2(G22gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n627_), .B2(new_n652_), .ZN(G1327gat));
  NAND2_X1  g452(.A1(new_n613_), .A2(new_n616_), .ZN(new_n654_));
  AND4_X1   g453(.A1(KEYINPUT98), .A2(new_n654_), .A3(new_n583_), .A4(new_n488_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT98), .B1(new_n617_), .B2(new_n488_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n622_), .A2(new_n625_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n423_), .A2(new_n425_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n451_), .A2(new_n206_), .A3(new_n452_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n257_), .A2(KEYINPUT33), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n456_), .B1(new_n455_), .B2(new_n256_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n660_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n440_), .A2(new_n442_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT93), .B1(new_n414_), .B2(new_n437_), .ZN(new_n665_));
  AOI211_X1 g464(.A(new_n445_), .B(new_n438_), .C1(new_n407_), .C2(new_n413_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n250_), .A2(new_n251_), .A3(new_n206_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n256_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n668_));
  OAI22_X1  g467(.A1(new_n665_), .A2(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  OAI22_X1  g468(.A1(new_n659_), .A2(new_n663_), .B1(new_n664_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n373_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT43), .B(new_n658_), .C1(new_n672_), .C2(new_n436_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  INV_X1    g473(.A(new_n658_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n460_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n657_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n657_), .B(KEYINPUT44), .C1(new_n673_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n619_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n617_), .A2(new_n488_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n460_), .A3(new_n562_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n684_), .A2(G29gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n682_), .B1(new_n619_), .B2(new_n685_), .ZN(G1328gat));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n679_), .A2(new_n636_), .A3(new_n680_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n679_), .A2(KEYINPUT99), .A3(new_n636_), .A4(new_n680_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(G36gat), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n684_), .A2(G36gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n636_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698_));
  INV_X1    g497(.A(new_n636_), .ZN(new_n699_));
  NOR4_X1   g498(.A1(new_n684_), .A2(KEYINPUT100), .A3(G36gat), .A4(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(new_n698_), .A3(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT45), .B1(new_n696_), .B2(new_n700_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n687_), .B(new_n688_), .C1(new_n693_), .C2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n687_), .A2(new_n688_), .ZN(new_n707_));
  AND4_X1   g506(.A1(new_n706_), .A2(new_n693_), .A3(new_n707_), .A4(new_n704_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1329gat));
  OAI21_X1  g508(.A(new_n491_), .B1(new_n684_), .B2(new_n644_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n326_), .A2(G43gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n681_), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g512(.A(G50gat), .B1(new_n681_), .B2(new_n649_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n370_), .A2(new_n489_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT102), .Z(new_n716_));
  OAI21_X1  g515(.A(new_n714_), .B1(new_n684_), .B2(new_n716_), .ZN(G1331gat));
  INV_X1    g516(.A(new_n654_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n626_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n584_), .B1(new_n719_), .B2(KEYINPUT103), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n461_), .B(new_n720_), .C1(KEYINPUT103), .C2(new_n719_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n258_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n654_), .A2(new_n583_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n563_), .A2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT104), .Z(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(KEYINPUT105), .A2(G57gat), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G57gat), .B1(new_n619_), .B2(KEYINPUT105), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n722_), .B1(new_n728_), .B2(new_n729_), .ZN(G1332gat));
  INV_X1    g529(.A(G64gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n721_), .A2(new_n731_), .A3(new_n636_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n725_), .A2(new_n636_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(G64gat), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT48), .B(new_n731_), .C1(new_n725_), .C2(new_n636_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n721_), .A2(new_n738_), .A3(new_n326_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT49), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n725_), .A2(new_n326_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(G71gat), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT49), .B(new_n738_), .C1(new_n725_), .C2(new_n326_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(G1334gat));
  INV_X1    g543(.A(G78gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n721_), .A2(new_n745_), .A3(new_n370_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n725_), .A2(new_n370_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(G78gat), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT50), .B(new_n745_), .C1(new_n725_), .C2(new_n370_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1335gat));
  OAI211_X1 g550(.A(new_n488_), .B(new_n723_), .C1(new_n673_), .C2(new_n676_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n619_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n723_), .A2(new_n488_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n461_), .A2(new_n754_), .A3(new_n561_), .ZN(new_n755_));
  INV_X1    g554(.A(G85gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n258_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n753_), .A2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT106), .ZN(G1336gat));
  AOI21_X1  g558(.A(G92gat), .B1(new_n755_), .B2(new_n636_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n752_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n636_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT107), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n760_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT108), .Z(G1337gat));
  OAI21_X1  g564(.A(G99gat), .B1(new_n752_), .B2(new_n644_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n644_), .A2(new_n528_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n755_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g569(.A1(new_n752_), .A2(new_n649_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT109), .B1(new_n771_), .B2(new_n507_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(G106gat), .C1(new_n752_), .C2(new_n649_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n774_), .A3(KEYINPUT52), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n755_), .A2(new_n507_), .A3(new_n370_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT109), .B(new_n777_), .C1(new_n771_), .C2(new_n507_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(G1339gat));
  XOR2_X1   g580(.A(KEYINPUT114), .B(G113gat), .Z(new_n782_));
  NAND2_X1  g581(.A1(new_n583_), .A2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT115), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT55), .B1(new_n597_), .B2(new_n600_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n596_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(G230gat), .A3(G233gat), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n598_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n607_), .B1(new_n785_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT56), .B(new_n607_), .C1(new_n785_), .C2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n564_), .A2(new_n571_), .A3(new_n568_), .A4(new_n569_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n565_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n579_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n582_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT112), .B1(new_n615_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n798_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n612_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n799_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n794_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n794_), .A2(new_n803_), .A3(KEYINPUT58), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n675_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n612_), .A2(new_n583_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n798_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n561_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT57), .B(new_n561_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n808_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n488_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n626_), .A2(new_n584_), .A3(new_n654_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n819_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n626_), .A2(new_n654_), .A3(new_n584_), .A4(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n370_), .B1(new_n817_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n699_), .A2(new_n258_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n644_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT59), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n823_), .B1(new_n816_), .B2(new_n488_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  INV_X1    g629(.A(new_n827_), .ZN(new_n831_));
  NOR4_X1   g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n370_), .A4(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n784_), .B1(new_n828_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n817_), .A2(new_n824_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(new_n583_), .A3(new_n649_), .A4(new_n827_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n211_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n835_), .B2(new_n211_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n833_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n833_), .B(KEYINPUT116), .C1(new_n837_), .C2(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1340gat));
  OAI21_X1  g642(.A(new_n718_), .B1(new_n828_), .B2(new_n832_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT117), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(new_n718_), .C1(new_n828_), .C2(new_n832_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(G120gat), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n834_), .A2(new_n649_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n831_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n215_), .B1(new_n654_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n850_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n215_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n852_), .ZN(G1341gat));
  INV_X1    g652(.A(new_n488_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G127gat), .B1(new_n850_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n828_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n832_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n488_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n855_), .B1(new_n858_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g658(.A(G134gat), .B1(new_n850_), .B2(new_n562_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT118), .B(G134gat), .Z(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n862_), .B2(new_n675_), .ZN(G1343gat));
  NOR3_X1   g662(.A1(new_n829_), .A2(new_n649_), .A3(new_n326_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n826_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n583_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n718_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g670(.A1(new_n866_), .A2(new_n488_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT61), .B(G155gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  NOR3_X1   g673(.A1(new_n866_), .A2(new_n553_), .A3(new_n658_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n553_), .B1(new_n866_), .B2(new_n561_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT119), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n878_), .B(new_n553_), .C1(new_n866_), .C2(new_n561_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n877_), .B2(new_n879_), .ZN(G1347gat));
  NAND3_X1  g679(.A1(new_n636_), .A2(new_n619_), .A3(new_n326_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT120), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n849_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n583_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G169gat), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n884_), .A2(G169gat), .A3(new_n886_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n383_), .A2(new_n389_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n888_), .B(new_n889_), .C1(new_n890_), .C2(new_n884_), .ZN(G1348gat));
  NAND2_X1  g690(.A1(new_n883_), .A2(new_n718_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g692(.A1(new_n883_), .A2(new_n854_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(G183gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n284_), .B1(KEYINPUT122), .B2(G183gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n894_), .B2(new_n897_), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n883_), .A2(new_n399_), .A3(new_n562_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n849_), .A2(new_n658_), .A3(new_n882_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n267_), .ZN(G1351gat));
  NAND3_X1  g700(.A1(new_n644_), .A2(new_n619_), .A3(new_n370_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n699_), .B1(new_n903_), .B2(KEYINPUT123), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n903_), .A2(KEYINPUT123), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n834_), .A2(new_n583_), .A3(new_n904_), .A4(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  OR3_X1    g706(.A1(new_n906_), .A2(new_n907_), .A3(KEYINPUT125), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT125), .B1(new_n906_), .B2(new_n907_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n906_), .A2(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(G197gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n908_), .A2(G197gat), .A3(new_n911_), .A4(new_n909_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1352gat));
  NAND3_X1  g714(.A1(new_n834_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n654_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(G204gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n917_), .B(new_n919_), .ZN(G1353gat));
  NAND4_X1  g719(.A1(new_n834_), .A2(new_n854_), .A3(new_n904_), .A4(new_n905_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n922_));
  INV_X1    g721(.A(G211gat), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  OR3_X1    g723(.A1(new_n921_), .A2(KEYINPUT127), .A3(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT127), .B1(new_n921_), .B2(new_n924_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n922_), .A2(new_n923_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n925_), .A2(new_n922_), .A3(new_n923_), .A4(new_n926_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1354gat));
  NOR2_X1   g730(.A1(new_n916_), .A2(new_n561_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(G218gat), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n916_), .A2(new_n658_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(G218gat), .B2(new_n934_), .ZN(G1355gat));
endmodule


