//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n940_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n972_, new_n973_, new_n974_, new_n976_, new_n977_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n984_, new_n985_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT17), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G155gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT16), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G183gat), .B(G211gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G64gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G57gat), .ZN(new_n209_));
  INV_X1    g008(.A(G57gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G64gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT11), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT69), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G57gat), .B(G64gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT11), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n210_), .A2(G64gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n208_), .A2(G57gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(G71gat), .A2(G78gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G71gat), .A2(G78gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT68), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT11), .B1(new_n209_), .B2(new_n211_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G71gat), .B(G78gat), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n217_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n227_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n224_), .B(KEYINPUT68), .C1(new_n214_), .C2(KEYINPUT11), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n213_), .A4(new_n216_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G1gat), .B(G8gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT73), .B(G15gat), .ZN(new_n237_));
  INV_X1    g036(.A(G22gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(G22gat), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G8gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n236_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n245_), .ZN(new_n247_));
  AOI211_X1 g046(.A(new_n235_), .B(new_n247_), .C1(new_n239_), .C2(new_n242_), .ZN(new_n248_));
  INV_X1    g047(.A(G231gat), .ZN(new_n249_));
  INV_X1    g048(.A(G233gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n246_), .A2(new_n248_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n242_), .ZN(new_n254_));
  AOI21_X1  g053(.A(G22gat), .B1(new_n240_), .B2(new_n241_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n245_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n235_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n243_), .A2(new_n236_), .A3(new_n245_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n253_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n234_), .B1(new_n252_), .B2(new_n259_), .ZN(new_n260_));
  AND4_X1   g059(.A1(new_n231_), .A2(new_n232_), .A3(new_n213_), .A4(new_n216_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n231_), .A2(new_n232_), .B1(new_n213_), .B2(new_n216_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n258_), .A3(new_n253_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n251_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n207_), .B1(new_n260_), .B2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT74), .B1(new_n260_), .B2(new_n266_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n207_), .ZN(new_n269_));
  OAI22_X1  g068(.A1(new_n203_), .A2(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n271_));
  INV_X1    g070(.A(new_n266_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(KEYINPUT17), .A3(new_n207_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT100), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G211gat), .B(G218gat), .Z(new_n281_));
  OR2_X1    g080(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n282_));
  INV_X1    g081(.A(G204gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(G197gat), .B2(G204gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n281_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G197gat), .A2(G204gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n288_), .B1(KEYINPUT21), .B2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT21), .A3(new_n281_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G183gat), .ZN(new_n300_));
  INV_X1    g099(.A(G190gat), .ZN(new_n301_));
  OAI211_X1 g100(.A(KEYINPUT83), .B(KEYINPUT23), .C1(new_n300_), .C2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT23), .B1(new_n300_), .B2(new_n301_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(G183gat), .A3(G190gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT83), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n299_), .A2(new_n302_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n301_), .A2(KEYINPUT26), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n301_), .A2(KEYINPUT26), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT95), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT26), .B(G190gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT95), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT25), .B(G183gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT97), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT24), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n296_), .B1(new_n320_), .B2(KEYINPUT96), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(KEYINPUT96), .B2(new_n320_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n317_), .A2(new_n318_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n318_), .B1(new_n317_), .B2(new_n322_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n309_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n303_), .A2(new_n305_), .A3(KEYINPUT81), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n327_), .A2(new_n304_), .A3(G183gat), .A4(G190gat), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(G183gat), .B2(G190gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n319_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT22), .B(G169gat), .ZN(new_n332_));
  INV_X1    g131(.A(G176gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n295_), .B1(new_n325_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT82), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT22), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n333_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT82), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(G169gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n307_), .B(new_n302_), .C1(G183gat), .C2(G190gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT24), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(G169gat), .B2(G176gat), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n316_), .A2(new_n313_), .B1(new_n346_), .B2(new_n297_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n329_), .B1(KEYINPUT80), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n316_), .A2(new_n313_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n297_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n299_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n344_), .B1(new_n348_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT20), .B1(new_n354_), .B2(new_n294_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n280_), .B1(new_n336_), .B2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT18), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n325_), .A2(new_n295_), .A3(new_n335_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n354_), .B2(new_n294_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n280_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n356_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT27), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n365_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n317_), .A2(new_n322_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT97), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n317_), .A2(new_n318_), .A3(new_n322_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n308_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n335_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n294_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n326_), .A2(new_n328_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n298_), .B1(new_n347_), .B2(KEYINPUT80), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n378_), .A2(new_n379_), .B1(new_n343_), .B2(new_n342_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n363_), .B1(new_n295_), .B2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n365_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n361_), .B1(new_n370_), .B2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n368_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n356_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n361_), .B1(new_n356_), .B2(new_n366_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT99), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n365_), .B1(new_n376_), .B2(new_n381_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n360_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n367_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(KEYINPUT99), .A3(new_n385_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n384_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  INV_X1    g199(.A(G155gat), .ZN(new_n401_));
  INV_X1    g200(.A(G162gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G141gat), .A2(G148gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT2), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT87), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n414_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417_));
  INV_X1    g216(.A(G141gat), .ZN(new_n418_));
  INV_X1    g217(.A(G148gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n411_), .A2(new_n416_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n406_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n411_), .A2(new_n416_), .A3(KEYINPUT88), .A4(new_n420_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n404_), .A2(KEYINPUT86), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT1), .B1(new_n401_), .B2(new_n402_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT1), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(G155gat), .A3(G162gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n403_), .A2(KEYINPUT86), .A3(new_n427_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n418_), .A2(new_n419_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n430_), .A2(new_n407_), .A3(new_n431_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n423_), .A2(new_n424_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G127gat), .B(G134gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT84), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G113gat), .B(G120gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n435_), .B(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n435_), .B(new_n436_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n413_), .A2(new_n415_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n420_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n422_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(new_n424_), .A3(new_n405_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n432_), .A2(new_n429_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n440_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G225gat), .A2(G233gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n439_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n439_), .A2(new_n447_), .A3(KEYINPUT4), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n440_), .A2(new_n446_), .A3(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n448_), .B(KEYINPUT98), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n400_), .B(new_n449_), .C1(new_n450_), .C2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n439_), .A2(new_n447_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n452_), .B(new_n453_), .C1(new_n457_), .C2(new_n451_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n400_), .B1(new_n458_), .B2(new_n449_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G228gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(new_n250_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT29), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n465_), .B2(new_n295_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT91), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT91), .B(new_n463_), .C1(new_n465_), .C2(new_n295_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n294_), .B1(new_n462_), .B2(new_n250_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n465_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n465_), .A2(KEYINPUT89), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G78gat), .B(G106gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT93), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n468_), .A2(new_n469_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n478_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n478_), .B(KEYINPUT92), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n470_), .A2(new_n484_), .A3(new_n476_), .ZN(new_n485_));
  OR3_X1    g284(.A1(new_n446_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT28), .B1(new_n446_), .B2(KEYINPUT29), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G22gat), .B(G50gat), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n479_), .A2(new_n483_), .A3(new_n485_), .A4(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n485_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n481_), .A2(new_n484_), .ZN(new_n494_));
  OAI22_X1  g293(.A1(new_n493_), .A2(new_n494_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n461_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n484_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n477_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n491_), .B1(new_n498_), .B2(new_n485_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n481_), .A2(new_n480_), .A3(new_n482_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n485_), .A2(new_n491_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n499_), .B1(new_n502_), .B2(new_n483_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n400_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n453_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n452_), .A2(new_n448_), .ZN(new_n506_));
  OAI221_X1 g305(.A(new_n504_), .B1(new_n457_), .B2(new_n505_), .C1(new_n450_), .C2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n393_), .A2(new_n507_), .A3(new_n367_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT33), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n455_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n458_), .A2(KEYINPUT33), .A3(new_n400_), .A4(new_n449_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n361_), .A2(KEYINPUT32), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n356_), .A2(new_n366_), .A3(new_n513_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n336_), .A2(new_n355_), .A3(new_n280_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(new_n369_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n514_), .B1(new_n516_), .B2(new_n513_), .ZN(new_n517_));
  OAI22_X1  g316(.A1(new_n508_), .A2(new_n512_), .B1(new_n460_), .B2(new_n517_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n396_), .A2(new_n496_), .B1(new_n503_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n440_), .B(KEYINPUT31), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G71gat), .B(G99gat), .ZN(new_n521_));
  INV_X1    g320(.A(G43gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n380_), .B(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G227gat), .A2(G233gat), .ZN(new_n525_));
  INV_X1    g324(.A(G15gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT30), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n524_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n520_), .B1(new_n530_), .B2(KEYINPUT85), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT85), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n529_), .A2(new_n532_), .A3(new_n520_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n277_), .B1(new_n519_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n518_), .A2(new_n495_), .A3(new_n492_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n492_), .A2(new_n495_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n460_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT99), .B1(new_n394_), .B2(new_n385_), .ZN(new_n542_));
  AOI211_X1 g341(.A(new_n389_), .B(KEYINPUT27), .C1(new_n393_), .C2(new_n367_), .ZN(new_n543_));
  OAI22_X1  g342(.A1(new_n542_), .A2(new_n543_), .B1(new_n383_), .B2(new_n368_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n539_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(KEYINPUT100), .A3(new_n536_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n536_), .A2(new_n461_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT101), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n396_), .A2(new_n548_), .ZN(new_n549_));
  AOI211_X1 g348(.A(KEYINPUT101), .B(new_n384_), .C1(new_n390_), .C2(new_n395_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n547_), .B(new_n503_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n538_), .A2(new_n546_), .A3(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G85gat), .B(G92gat), .Z(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT9), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT65), .B(G92gat), .ZN(new_n555_));
  INV_X1    g354(.A(G85gat), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(KEYINPUT9), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT6), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT6), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(G99gat), .A3(G106gat), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n555_), .A2(new_n557_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT10), .B(G99gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(G106gat), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT64), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT64), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n563_), .A2(new_n567_), .A3(G106gat), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n554_), .B(new_n562_), .C1(new_n566_), .C2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT8), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n559_), .A2(new_n561_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT67), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT67), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n559_), .A2(new_n561_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n575_));
  INV_X1    g374(.A(G99gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n565_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n572_), .A2(new_n574_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n570_), .B1(new_n580_), .B2(new_n553_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n570_), .A2(KEYINPUT66), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n570_), .A2(KEYINPUT66), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n553_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n571_), .B2(new_n579_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n569_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G29gat), .B(G36gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G43gat), .B(G50gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT15), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n587_), .A2(new_n588_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n587_), .A2(new_n588_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(KEYINPUT15), .A3(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n586_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n579_), .A2(new_n571_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n597_), .A2(new_n553_), .A3(new_n582_), .A4(new_n583_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n553_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n573_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n577_), .A2(new_n578_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n599_), .B1(new_n602_), .B2(new_n574_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n598_), .B1(new_n603_), .B2(new_n570_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n569_), .A3(new_n589_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT34), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n596_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n608_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n596_), .A2(new_n605_), .A3(new_n612_), .A4(new_n609_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G134gat), .B(G162gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(KEYINPUT36), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n617_), .B(KEYINPUT36), .Z(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n614_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n586_), .A2(new_n263_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n234_), .B1(new_n604_), .B2(new_n569_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT12), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT12), .B1(new_n586_), .B2(new_n263_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n629_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(G120gat), .B(G148gat), .Z(new_n636_));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n635_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n640_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n632_), .A2(new_n634_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT13), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n641_), .A2(KEYINPUT13), .A3(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n591_), .B(new_n594_), .C1(new_n246_), .C2(new_n248_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n257_), .A2(new_n258_), .A3(new_n589_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(KEYINPUT77), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT77), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n257_), .A2(new_n258_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n595_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n650_), .B1(new_n653_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT76), .ZN(new_n658_));
  INV_X1    g457(.A(new_n589_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n659_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n660_));
  AOI211_X1 g459(.A(new_n658_), .B(new_n649_), .C1(new_n660_), .C2(new_n652_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n652_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT76), .B1(new_n662_), .B2(new_n650_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n657_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(G113gat), .B(G141gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(G169gat), .B(G197gat), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n665_), .B(new_n666_), .Z(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT78), .B1(new_n664_), .B2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n663_), .A2(new_n661_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n653_), .A2(new_n656_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n649_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT78), .ZN(new_n673_));
  INV_X1    g472(.A(new_n667_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT79), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n664_), .A2(new_n676_), .A3(new_n667_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n669_), .A2(new_n671_), .A3(new_n667_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT79), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n668_), .A2(new_n675_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n648_), .A2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT102), .ZN(new_n682_));
  AND4_X1   g481(.A1(new_n276_), .A2(new_n552_), .A3(new_n625_), .A4(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n202_), .B1(new_n683_), .B2(new_n461_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n552_), .A2(new_n681_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n619_), .B(new_n686_), .C1(new_n614_), .C2(new_n622_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n270_), .A2(new_n275_), .A3(KEYINPUT75), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT75), .B1(new_n270_), .B2(new_n275_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n691_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n685_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n202_), .A3(new_n461_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT38), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n684_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n699_), .B1(new_n698_), .B2(new_n697_), .ZN(G1324gat));
  NOR2_X1   g499(.A1(new_n549_), .A2(new_n550_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n683_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G8gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT39), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n696_), .A2(new_n244_), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(G1325gat));
  AOI21_X1  g507(.A(new_n526_), .B1(new_n683_), .B2(new_n537_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT41), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n696_), .A2(new_n526_), .A3(new_n537_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1326gat));
  NAND2_X1  g511(.A1(new_n683_), .A2(new_n540_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G22gat), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT42), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n696_), .A2(new_n238_), .A3(new_n540_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT103), .ZN(G1327gat));
  OR2_X1    g517(.A1(new_n692_), .A2(new_n693_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n625_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n685_), .A2(new_n720_), .ZN(new_n721_));
  OR3_X1    g520(.A1(new_n721_), .A2(G29gat), .A3(new_n460_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n682_), .A2(new_n694_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n552_), .A2(new_n724_), .A3(new_n691_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n552_), .B2(new_n691_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n723_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT44), .B(new_n723_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n461_), .A3(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n729_), .A2(KEYINPUT104), .A3(new_n461_), .A4(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G29gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n722_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT105), .B(new_n722_), .C1(new_n733_), .C2(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1328gat));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n701_), .A2(KEYINPUT106), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n701_), .A2(KEYINPUT106), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n721_), .A2(G36gat), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n729_), .A2(new_n701_), .A3(new_n730_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G36gat), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n741_), .B(new_n742_), .C1(new_n749_), .C2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n741_), .A2(new_n742_), .ZN(new_n754_));
  AND4_X1   g553(.A1(new_n753_), .A2(new_n749_), .A3(new_n751_), .A4(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1329gat));
  NAND3_X1  g555(.A1(new_n685_), .A2(new_n537_), .A3(new_n720_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT109), .A3(new_n522_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT109), .B1(new_n757_), .B2(new_n522_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n536_), .A2(new_n522_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n729_), .A2(new_n730_), .A3(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n729_), .A2(KEYINPUT108), .A3(new_n730_), .A4(new_n761_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n760_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n766_), .B(new_n768_), .ZN(G1330gat));
  AND2_X1   g568(.A1(new_n729_), .A2(new_n730_), .ZN(new_n770_));
  INV_X1    g569(.A(G50gat), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n503_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n685_), .A2(new_n540_), .A3(new_n720_), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n770_), .A2(new_n772_), .B1(new_n771_), .B2(new_n773_), .ZN(G1331gat));
  AND2_X1   g573(.A1(new_n646_), .A2(new_n647_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n668_), .A2(new_n675_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n677_), .A2(new_n679_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n775_), .A2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n552_), .A2(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n780_), .A2(new_n719_), .A3(new_n625_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n210_), .B1(new_n781_), .B2(new_n461_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n780_), .A2(new_n695_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n460_), .A2(G57gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT111), .Z(G1332gat));
  AOI21_X1  g585(.A(new_n208_), .B1(new_n781_), .B2(new_n745_), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT48), .Z(new_n788_));
  NAND3_X1  g587(.A1(new_n783_), .A2(new_n208_), .A3(new_n745_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1333gat));
  INV_X1    g589(.A(G71gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n781_), .B2(new_n537_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT49), .Z(new_n793_));
  NAND3_X1  g592(.A1(new_n783_), .A2(new_n791_), .A3(new_n537_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(G1334gat));
  INV_X1    g594(.A(G78gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(new_n781_), .B2(new_n540_), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT50), .Z(new_n798_));
  NAND3_X1  g597(.A1(new_n783_), .A2(new_n796_), .A3(new_n540_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1335gat));
  NAND2_X1  g599(.A1(new_n780_), .A2(new_n720_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G85gat), .B1(new_n803_), .B2(new_n461_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n725_), .A2(new_n726_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n779_), .A2(new_n694_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n460_), .A2(new_n556_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT113), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n804_), .B1(new_n807_), .B2(new_n809_), .ZN(G1336gat));
  AOI21_X1  g609(.A(G92gat), .B1(new_n803_), .B2(new_n701_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n745_), .A2(new_n555_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n807_), .B2(new_n812_), .ZN(G1337gat));
  NOR2_X1   g612(.A1(new_n536_), .A2(new_n563_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n803_), .A2(new_n814_), .B1(new_n815_), .B2(KEYINPUT51), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n807_), .A2(new_n537_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G99gat), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n815_), .A2(KEYINPUT51), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1338gat));
  NAND3_X1  g620(.A1(new_n803_), .A2(new_n565_), .A3(new_n540_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n807_), .A2(new_n540_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(G106gat), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT52), .B(new_n565_), .C1(new_n807_), .C2(new_n540_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n822_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT53), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n829_), .B(new_n822_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1339gat));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  NOR4_X1   g631(.A1(new_n701_), .A2(new_n536_), .A3(new_n460_), .A4(new_n540_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n778_), .A2(new_n643_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT12), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n586_), .A2(new_n263_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n604_), .A2(new_n234_), .A3(new_n569_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841_));
  NOR4_X1   g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n633_), .A4(new_n630_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n629_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n840_), .A2(new_n633_), .A3(new_n630_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT116), .B1(new_n845_), .B2(KEYINPUT55), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n632_), .A2(new_n847_), .A3(new_n841_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n844_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n640_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(KEYINPUT56), .A3(new_n640_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n836_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n650_), .B1(new_n660_), .B2(new_n652_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n667_), .B(new_n855_), .C1(new_n670_), .C2(new_n650_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n644_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n625_), .B1(new_n854_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n643_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n849_), .A2(KEYINPUT56), .A3(new_n640_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT56), .B1(new_n849_), .B2(new_n640_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n690_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n864_), .B(KEYINPUT58), .C1(new_n865_), .C2(new_n866_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n861_), .A2(new_n860_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n862_), .B1(new_n871_), .B2(KEYINPUT117), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n860_), .A2(new_n861_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n869_), .A2(new_n870_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n873_), .A2(KEYINPUT117), .A3(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n694_), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n778_), .A2(new_n694_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n775_), .A2(KEYINPUT115), .A3(new_n877_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n719_), .A2(new_n646_), .A3(new_n680_), .A4(new_n647_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n881_), .A3(new_n690_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT54), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n878_), .A2(new_n881_), .A3(new_n884_), .A4(new_n690_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n835_), .B1(new_n876_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n276_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n873_), .A2(new_n874_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n860_), .A2(new_n861_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n887_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n834_), .B1(new_n893_), .B2(new_n833_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n832_), .B1(new_n888_), .B2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n871_), .A2(new_n862_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n886_), .B1(new_n896_), .B2(new_n889_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n833_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT59), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n890_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n871_), .A2(KEYINPUT117), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n902_), .A3(new_n862_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n886_), .B1(new_n903_), .B2(new_n694_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n899_), .B(KEYINPUT118), .C1(new_n904_), .C2(new_n835_), .ZN(new_n905_));
  INV_X1    g704(.A(G113gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n680_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n895_), .A2(new_n905_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n893_), .A2(new_n833_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n909_), .B2(new_n680_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n908_), .A2(KEYINPUT119), .A3(new_n910_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1340gat));
  OAI21_X1  g714(.A(new_n899_), .B1(new_n904_), .B2(new_n835_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G120gat), .B1(new_n916_), .B2(new_n775_), .ZN(new_n917_));
  INV_X1    g716(.A(G120gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n775_), .B2(KEYINPUT60), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n919_), .B1(KEYINPUT60), .B2(new_n918_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n917_), .B1(new_n909_), .B2(new_n920_), .ZN(G1341gat));
  XOR2_X1   g720(.A(KEYINPUT120), .B(G127gat), .Z(new_n922_));
  NOR2_X1   g721(.A1(new_n889_), .A2(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n895_), .A2(new_n905_), .A3(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(G127gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n909_), .B2(new_n694_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT121), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n924_), .A2(new_n929_), .A3(new_n926_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1342gat));
  NAND3_X1  g730(.A1(new_n895_), .A2(new_n905_), .A3(new_n691_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(G134gat), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n625_), .A2(G134gat), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n909_), .B2(new_n934_), .ZN(G1343gat));
  NOR2_X1   g734(.A1(new_n897_), .A2(new_n537_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n936_), .A2(new_n461_), .A3(new_n540_), .A4(new_n746_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n680_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n418_), .ZN(G1344gat));
  NOR2_X1   g738(.A1(new_n937_), .A2(new_n775_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(new_n419_), .ZN(G1345gat));
  NOR2_X1   g740(.A1(new_n937_), .A2(new_n694_), .ZN(new_n942_));
  XOR2_X1   g741(.A(KEYINPUT61), .B(G155gat), .Z(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1346gat));
  NOR3_X1   g743(.A1(new_n937_), .A2(new_n402_), .A3(new_n690_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n402_), .B1(new_n937_), .B2(new_n625_), .ZN(new_n946_));
  OR2_X1    g745(.A1(new_n946_), .A2(KEYINPUT122), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(KEYINPUT122), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n945_), .B1(new_n947_), .B2(new_n948_), .ZN(G1347gat));
  NAND2_X1  g748(.A1(new_n876_), .A2(new_n887_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n745_), .A2(new_n547_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(KEYINPUT123), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n745_), .A2(new_n953_), .A3(new_n547_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n540_), .B1(new_n952_), .B2(new_n954_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n950_), .A2(new_n778_), .A3(new_n955_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(G169gat), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n956_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n959_), .A2(KEYINPUT62), .A3(new_n960_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n957_), .A2(new_n958_), .A3(new_n962_), .ZN(new_n963_));
  AND2_X1   g762(.A1(new_n950_), .A2(new_n955_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n964_), .A2(new_n778_), .A3(new_n332_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n961_), .A2(new_n963_), .A3(new_n965_), .ZN(G1348gat));
  AOI21_X1  g765(.A(G176gat), .B1(new_n964_), .B2(new_n648_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n893_), .A2(new_n503_), .ZN(new_n968_));
  INV_X1    g767(.A(new_n968_), .ZN(new_n969_));
  AOI211_X1 g768(.A(new_n333_), .B(new_n775_), .C1(new_n952_), .C2(new_n954_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n967_), .B1(new_n969_), .B2(new_n970_), .ZN(G1349gat));
  AOI21_X1  g770(.A(new_n694_), .B1(new_n952_), .B2(new_n954_), .ZN(new_n972_));
  AOI21_X1  g771(.A(G183gat), .B1(new_n969_), .B2(new_n972_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n889_), .A2(new_n316_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n973_), .B1(new_n964_), .B2(new_n974_), .ZN(G1350gat));
  NAND4_X1  g774(.A1(new_n964_), .A2(new_n624_), .A3(new_n312_), .A4(new_n315_), .ZN(new_n976_));
  AND2_X1   g775(.A1(new_n964_), .A2(new_n691_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n977_), .B2(new_n301_), .ZN(G1351gat));
  NOR2_X1   g777(.A1(new_n746_), .A2(new_n541_), .ZN(new_n979_));
  AND2_X1   g778(.A1(new_n936_), .A2(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n980_), .A2(new_n778_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n983_));
  OAI211_X1 g782(.A(new_n980_), .B(new_n648_), .C1(new_n983_), .C2(new_n283_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n983_), .A2(new_n283_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n984_), .B(new_n985_), .ZN(G1353gat));
  NAND2_X1  g785(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n987_));
  OR3_X1    g786(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988_));
  NAND4_X1  g787(.A1(new_n980_), .A2(new_n276_), .A3(new_n987_), .A4(new_n988_), .ZN(new_n989_));
  OAI21_X1  g788(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n990_));
  XOR2_X1   g789(.A(new_n989_), .B(new_n990_), .Z(G1354gat));
  INV_X1    g790(.A(G218gat), .ZN(new_n992_));
  NAND3_X1  g791(.A1(new_n980_), .A2(new_n992_), .A3(new_n624_), .ZN(new_n993_));
  AND3_X1   g792(.A1(new_n936_), .A2(new_n691_), .A3(new_n979_), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n993_), .B1(new_n992_), .B2(new_n994_), .ZN(new_n995_));
  NAND2_X1  g794(.A1(new_n995_), .A2(KEYINPUT127), .ZN(new_n996_));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n997_));
  OAI211_X1 g796(.A(new_n993_), .B(new_n997_), .C1(new_n992_), .C2(new_n994_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n996_), .A2(new_n998_), .ZN(G1355gat));
endmodule


