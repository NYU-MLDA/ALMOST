//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206_));
  NOR3_X1   g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n207_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT10), .B(G99gat), .Z(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n204_), .A2(new_n206_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n213_), .A2(new_n214_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  AND3_X1   g018(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  INV_X1    g022(.A(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT9), .A3(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n227_), .A3(new_n218_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT10), .B(G99gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(G106gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(G99gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n216_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n235_), .A2(new_n210_), .A3(new_n211_), .A4(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n204_), .A2(new_n205_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n232_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n237_), .A2(new_n232_), .A3(new_n238_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n219_), .B(new_n231_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G57gat), .ZN(new_n242_));
  INV_X1    g041(.A(G64gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G57gat), .A2(G64gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT11), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G71gat), .B(G78gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n244_), .A2(new_n250_), .A3(new_n245_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT11), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT12), .B1(new_n241_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n241_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n256_), .A2(KEYINPUT67), .B1(new_n257_), .B2(new_n254_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT67), .B1(new_n241_), .B2(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n219_), .A2(new_n231_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n240_), .A2(new_n239_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT65), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n239_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n237_), .A2(new_n232_), .A3(new_n238_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(new_n219_), .A4(new_n231_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n254_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n252_), .A2(KEYINPUT66), .A3(new_n253_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n259_), .B1(new_n268_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT12), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n203_), .B(new_n258_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n257_), .A2(new_n254_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n241_), .A2(new_n255_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(G230gat), .A3(G233gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(G120gat), .B(G148gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G176gat), .B(G204gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n276_), .A2(new_n280_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n202_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n276_), .A2(new_n280_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n285_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n276_), .A2(new_n280_), .A3(new_n286_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT13), .A3(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G22gat), .ZN(new_n295_));
  INV_X1    g094(.A(G1gat), .ZN(new_n296_));
  INV_X1    g095(.A(G8gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT14), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G29gat), .A2(G36gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G43gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G29gat), .A2(G36gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n305_), .ZN(new_n307_));
  OAI21_X1  g106(.A(G43gat), .B1(new_n307_), .B2(new_n302_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n306_), .A2(new_n308_), .A3(G50gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(G50gat), .B1(new_n306_), .B2(new_n308_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n311_), .A2(KEYINPUT74), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(KEYINPUT74), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n301_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT15), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n309_), .A2(new_n310_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n306_), .A2(new_n308_), .ZN(new_n319_));
  INV_X1    g118(.A(G50gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n306_), .A2(new_n308_), .A3(G50gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT15), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n301_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n315_), .A2(new_n316_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n316_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n312_), .A2(new_n301_), .A3(new_n313_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n329_), .B2(new_n314_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G113gat), .B(G141gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G197gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT75), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G169gat), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n327_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n301_), .B(new_n254_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G231gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT72), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n339_), .B(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G127gat), .B(G155gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G183gat), .B(G211gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n342_), .B1(KEYINPUT17), .B2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n269_), .A3(KEYINPUT17), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n294_), .A2(new_n338_), .A3(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT71), .B(KEYINPUT37), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n324_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n241_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G232gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT34), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(KEYINPUT35), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n355_), .A2(new_n356_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n268_), .A2(new_n325_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT70), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(KEYINPUT35), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT69), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G190gat), .B(G218gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G134gat), .ZN(new_n368_));
  INV_X1    g167(.A(G162gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT36), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n356_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n359_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n361_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n365_), .B1(new_n355_), .B2(KEYINPUT70), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n366_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n370_), .A2(new_n371_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n366_), .B2(new_n377_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n354_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n375_), .A2(new_n376_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n375_), .A2(new_n376_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n379_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n366_), .A2(new_n377_), .A3(new_n372_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n353_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G169gat), .ZN(new_n389_));
  INV_X1    g188(.A(G176gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT22), .B(G169gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(new_n390_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(KEYINPUT23), .B2(new_n395_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n393_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n395_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(KEYINPUT23), .B2(new_n395_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT24), .B1(new_n389_), .B2(new_n390_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403_));
  MUX2_X1   g202(.A(new_n402_), .B(KEYINPUT24), .S(new_n403_), .Z(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT25), .B(G183gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n406_));
  INV_X1    g205(.A(G190gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(KEYINPUT26), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT26), .B(G190gat), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n405_), .B(new_n408_), .C1(new_n409_), .C2(new_n406_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n401_), .A2(new_n404_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n399_), .A2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n412_), .B(KEYINPUT30), .Z(new_n413_));
  OR2_X1    g212(.A1(new_n413_), .A2(new_n234_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n234_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G227gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G71gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G15gat), .B(G43gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n416_), .A2(new_n420_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G127gat), .B(G134gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G113gat), .B(G120gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT78), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n424_), .B(new_n426_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n429_), .B1(new_n430_), .B2(new_n428_), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n431_), .B(KEYINPUT31), .Z(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(KEYINPUT79), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n432_), .A2(KEYINPUT79), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n421_), .B(new_n423_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n421_), .ZN(new_n436_));
  OAI22_X1  g235(.A1(new_n436_), .A2(new_n422_), .B1(KEYINPUT79), .B2(new_n432_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT81), .A2(G228gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(KEYINPUT81), .A2(G228gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(G233gat), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G211gat), .B(G218gat), .Z(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT21), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G197gat), .B(G204gat), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT84), .B(KEYINPUT21), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n444_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n447_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(G197gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(G204gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n446_), .B1(new_n455_), .B2(KEYINPUT82), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(KEYINPUT83), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT83), .B1(new_n453_), .B2(new_n456_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n451_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n453_), .A2(new_n456_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT83), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n457_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT85), .B1(new_n466_), .B2(new_n451_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n449_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT29), .ZN(new_n469_));
  AND2_X1   g268(.A1(G155gat), .A2(G162gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G155gat), .A2(G162gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT1), .ZN(new_n473_));
  INV_X1    g272(.A(G141gat), .ZN(new_n474_));
  INV_X1    g273(.A(G148gat), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n472_), .A2(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n470_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OR3_X1    g277(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT2), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n479_), .A2(new_n481_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n472_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n469_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n443_), .B1(new_n468_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT80), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n478_), .A2(new_n489_), .A3(new_n485_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n443_), .B1(new_n492_), .B2(new_n469_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n460_), .A2(new_n461_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n466_), .A2(KEYINPUT85), .A3(new_n451_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n448_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G22gat), .B(G50gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT28), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n488_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n492_), .A2(new_n469_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G78gat), .B(G106gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  OAI21_X1  g303(.A(new_n499_), .B1(new_n488_), .B2(new_n497_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n504_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n505_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n507_), .B1(new_n508_), .B2(new_n500_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n412_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n512_), .B(new_n449_), .C1(new_n462_), .C2(new_n467_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n409_), .A2(new_n405_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n397_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n404_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n401_), .B1(G183gat), .B2(G190gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n393_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n513_), .B(KEYINPUT20), .C1(new_n496_), .C2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G226gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT19), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT18), .B(G64gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G92gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G8gat), .B(G36gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(KEYINPUT20), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n496_), .B2(new_n521_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n524_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n468_), .A2(new_n412_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n525_), .A2(new_n529_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n529_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n530_), .B1(new_n468_), .B2(new_n520_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n532_), .B1(new_n537_), .B2(new_n513_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT20), .B1(new_n468_), .B2(new_n520_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n532_), .B1(new_n496_), .B2(new_n512_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n536_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n535_), .A2(new_n542_), .A3(KEYINPUT86), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n525_), .A2(new_n534_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT86), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n536_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT0), .B(G57gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(G85gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(G1gat), .B(G29gat), .Z(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G225gat), .A2(G233gat), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n430_), .A2(KEYINPUT88), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n430_), .A2(KEYINPUT88), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n478_), .A2(new_n485_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(KEYINPUT80), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n478_), .A2(new_n489_), .A3(new_n485_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT87), .B1(new_n561_), .B2(new_n431_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n431_), .B(KEYINPUT87), .C1(new_n490_), .C2(new_n491_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(KEYINPUT4), .B(new_n558_), .C1(new_n562_), .C2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT89), .B(KEYINPUT4), .Z(new_n566_));
  NAND3_X1  g365(.A1(new_n561_), .A2(new_n431_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n553_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n431_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT87), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n557_), .B1(new_n571_), .B2(new_n563_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n553_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n552_), .B1(new_n568_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT90), .B(KEYINPUT33), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  OAI211_X1 g379(.A(KEYINPUT33), .B(new_n552_), .C1(new_n568_), .C2(new_n574_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT92), .ZN(new_n582_));
  AOI211_X1 g381(.A(new_n553_), .B(new_n557_), .C1(new_n571_), .C2(new_n563_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n582_), .B1(new_n583_), .B2(new_n552_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n572_), .A2(new_n573_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(KEYINPUT92), .A3(new_n551_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n565_), .A2(new_n553_), .A3(new_n567_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n584_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n581_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n575_), .A2(KEYINPUT91), .A3(new_n577_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n547_), .A2(new_n580_), .A3(new_n589_), .A4(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT94), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT93), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n533_), .B1(new_n531_), .B2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n539_), .A2(KEYINPUT93), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n592_), .B(new_n524_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n529_), .A2(KEYINPUT32), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n539_), .A2(KEYINPUT93), .B1(new_n468_), .B2(new_n412_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n531_), .A2(new_n593_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n532_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT94), .B1(new_n522_), .B2(new_n524_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n596_), .B(new_n597_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n568_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n574_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n551_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n575_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n602_), .B(new_n606_), .C1(new_n544_), .C2(new_n597_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n511_), .B1(new_n591_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n510_), .A2(new_n606_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n596_), .B(new_n536_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(KEYINPUT27), .A3(new_n535_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT27), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n543_), .A2(new_n546_), .A3(new_n612_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n609_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n439_), .B1(new_n608_), .B2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n606_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n611_), .A2(KEYINPUT95), .A3(new_n613_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT95), .B1(new_n611_), .B2(new_n613_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n510_), .B(new_n616_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  AOI211_X1 g418(.A(new_n352_), .B(new_n388_), .C1(new_n615_), .C2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n296_), .A3(new_n606_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT38), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n615_), .A2(new_n619_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n352_), .A2(KEYINPUT96), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n352_), .A2(KEYINPUT96), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n385_), .A2(new_n386_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n623_), .A2(new_n625_), .A3(new_n626_), .A4(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n606_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n622_), .A2(new_n631_), .ZN(G1324gat));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n617_), .A2(new_n618_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n633_), .B1(new_n629_), .B2(new_n635_), .ZN(new_n636_));
  AOI211_X1 g435(.A(new_n624_), .B(new_n627_), .C1(new_n615_), .C2(new_n619_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n637_), .A2(KEYINPUT97), .A3(new_n626_), .A4(new_n634_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(new_n638_), .A3(G8gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT98), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n636_), .A2(new_n638_), .A3(new_n641_), .A4(G8gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n620_), .A2(new_n297_), .A3(new_n634_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n640_), .A2(KEYINPUT39), .A3(new_n642_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n645_), .A2(new_n649_), .A3(new_n646_), .A4(new_n647_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n629_), .B2(new_n439_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT41), .Z(new_n655_));
  INV_X1    g454(.A(G15gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n620_), .A2(new_n656_), .A3(new_n438_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT100), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(G1326gat));
  OAI21_X1  g458(.A(G22gat), .B1(new_n629_), .B2(new_n510_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n620_), .A2(new_n662_), .A3(new_n511_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1327gat));
  AOI21_X1  g463(.A(new_n628_), .B1(new_n615_), .B2(new_n619_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n294_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n666_), .A2(new_n337_), .A3(new_n351_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n606_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n623_), .B2(new_n388_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n388_), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT43), .B(new_n672_), .C1(new_n615_), .C2(new_n619_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n667_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(G29gat), .ZN(new_n677_));
  OAI211_X1 g476(.A(KEYINPUT44), .B(new_n667_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(new_n606_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n669_), .B1(new_n677_), .B2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n668_), .A2(new_n681_), .A3(new_n634_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT45), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n672_), .B1(new_n615_), .B2(new_n619_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(new_n670_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT44), .B1(new_n686_), .B2(new_n667_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n678_), .A2(new_n634_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n684_), .B(G36gat), .C1(new_n687_), .C2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n676_), .A2(new_n634_), .A3(new_n678_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n684_), .B1(new_n691_), .B2(G36gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n683_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT46), .B(new_n683_), .C1(new_n690_), .C2(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1329gat));
  INV_X1    g496(.A(new_n668_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n304_), .B1(new_n698_), .B2(new_n439_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n676_), .A2(G43gat), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n678_), .A2(new_n438_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g502(.A1(new_n678_), .A2(new_n511_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G50gat), .B1(new_n687_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n511_), .A2(new_n320_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT102), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n698_), .B2(new_n707_), .ZN(G1331gat));
  NOR2_X1   g507(.A1(new_n294_), .A2(new_n338_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n623_), .A2(new_n709_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n382_), .A2(new_n351_), .A3(new_n387_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n606_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n710_), .A2(new_n351_), .A3(new_n628_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n715_), .A2(new_n242_), .A3(new_n630_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n715_), .B2(new_n635_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT103), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n720_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n713_), .A2(new_n243_), .A3(new_n634_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(G1333gat));
  OAI21_X1  g523(.A(G71gat), .B1(new_n715_), .B2(new_n439_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT49), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n439_), .A2(G71gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n712_), .B2(new_n727_), .ZN(G1334gat));
  OAI21_X1  g527(.A(G78gat), .B1(new_n715_), .B2(new_n510_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT50), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n510_), .A2(G78gat), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT104), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n712_), .B2(new_n732_), .ZN(G1335gat));
  INV_X1    g532(.A(new_n351_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n709_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n686_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737_), .B2(new_n630_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n665_), .A2(new_n736_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n223_), .A3(new_n606_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT105), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n740_), .B2(new_n634_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n686_), .A2(G92gat), .A3(new_n736_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n746_), .B2(new_n634_), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n737_), .B2(new_n439_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n740_), .A2(new_n215_), .A3(new_n438_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g550(.A(new_n511_), .B(new_n736_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G106gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT107), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n755_), .A3(G106gat), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT106), .B(KEYINPUT52), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n754_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n740_), .A2(new_n216_), .A3(new_n511_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n756_), .A2(new_n757_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(G1339gat));
  NAND3_X1  g562(.A1(new_n382_), .A2(new_n387_), .A3(new_n351_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n289_), .A2(new_n293_), .A3(new_n337_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(KEYINPUT109), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT109), .B1(new_n764_), .B2(new_n765_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n767_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n289_), .A2(new_n293_), .A3(new_n337_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n711_), .B2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT110), .B1(new_n776_), .B2(KEYINPUT54), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n766_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n773_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n272_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT12), .B1(new_n781_), .B2(new_n259_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n203_), .B1(new_n782_), .B2(new_n258_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n276_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n256_), .A2(KEYINPUT67), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n277_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n268_), .A2(new_n273_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n259_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n787_), .B1(new_n790_), .B2(KEYINPUT12), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(new_n203_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n276_), .B2(new_n784_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n785_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n285_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT56), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n798_), .A3(new_n285_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n797_), .A2(new_n338_), .A3(new_n292_), .A4(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n315_), .A2(new_n328_), .A3(new_n326_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n316_), .B1(new_n329_), .B2(new_n314_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n334_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n804_), .A2(new_n805_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n335_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n288_), .B2(new_n287_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n800_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n628_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(KEYINPUT57), .A3(new_n628_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n799_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n798_), .B1(new_n795_), .B2(new_n285_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n815_), .A2(new_n287_), .A3(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(KEYINPUT58), .A3(new_n808_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n797_), .A2(new_n292_), .A3(new_n808_), .A4(new_n799_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n821_), .A3(new_n388_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n813_), .A2(new_n814_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n780_), .B1(new_n823_), .B2(new_n734_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n510_), .B(new_n438_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n606_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT113), .B1(new_n825_), .B2(new_n630_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n824_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(new_n338_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n823_), .A2(new_n734_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n780_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n830_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n824_), .B2(KEYINPUT114), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n832_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n338_), .A2(G113gat), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT115), .Z(new_n846_));
  AOI21_X1  g645(.A(new_n833_), .B1(new_n844_), .B2(new_n846_), .ZN(G1340gat));
  AOI221_X4 g646(.A(new_n831_), .B1(KEYINPUT114), .B2(new_n840_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n842_), .A2(new_n832_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n666_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT116), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n844_), .A2(new_n852_), .A3(new_n666_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n851_), .A2(G120gat), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n294_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n832_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(G1341gat));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859_));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  AOI211_X1 g659(.A(new_n860_), .B(new_n734_), .C1(new_n841_), .C2(new_n843_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n837_), .B2(new_n734_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT117), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n864_), .B(new_n860_), .C1(new_n837_), .C2(new_n734_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n859_), .B1(new_n861_), .B2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n844_), .A2(G127gat), .A3(new_n351_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n868_), .A2(KEYINPUT118), .A3(new_n865_), .A4(new_n863_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(G1342gat));
  INV_X1    g669(.A(G134gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n837_), .B2(new_n628_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n872_), .A2(KEYINPUT119), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(KEYINPUT119), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n388_), .A2(G134gat), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT120), .Z(new_n876_));
  AOI22_X1  g675(.A1(new_n873_), .A2(new_n874_), .B1(new_n844_), .B2(new_n876_), .ZN(G1343gat));
  NOR2_X1   g676(.A1(new_n438_), .A2(new_n510_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n824_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n634_), .A2(new_n630_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n337_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n474_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n294_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n475_), .ZN(G1345gat));
  NOR2_X1   g685(.A1(new_n882_), .A2(new_n734_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT61), .B(G155gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  NOR3_X1   g688(.A1(new_n882_), .A2(new_n369_), .A3(new_n672_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n880_), .A2(new_n627_), .A3(new_n881_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n369_), .B2(new_n891_), .ZN(G1347gat));
  AOI21_X1  g691(.A(new_n635_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(new_n510_), .A3(new_n616_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n337_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n896_), .A2(KEYINPUT121), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(KEYINPUT121), .ZN(new_n898_));
  OR4_X1    g697(.A1(new_n389_), .A2(new_n895_), .A3(new_n897_), .A4(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n392_), .ZN(new_n900_));
  OAI211_X1 g699(.A(KEYINPUT121), .B(new_n896_), .C1(new_n895_), .C2(new_n389_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(G1348gat));
  NOR2_X1   g701(.A1(new_n894_), .A2(new_n294_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT122), .B(G176gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1349gat));
  NOR2_X1   g704(.A1(new_n894_), .A2(new_n734_), .ZN(new_n906_));
  MUX2_X1   g705(.A(G183gat), .B(new_n405_), .S(new_n906_), .Z(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n894_), .B2(new_n672_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n627_), .A2(new_n409_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n894_), .B2(new_n909_), .ZN(G1351gat));
  NOR2_X1   g709(.A1(new_n879_), .A2(new_n606_), .ZN(new_n911_));
  AOI21_X1  g710(.A(KEYINPUT57), .B1(new_n810_), .B2(new_n628_), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n812_), .B(new_n627_), .C1(new_n800_), .C2(new_n809_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n351_), .B1(new_n914_), .B2(new_n822_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n634_), .B(new_n911_), .C1(new_n915_), .C2(new_n780_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n836_), .A2(KEYINPUT123), .A3(new_n634_), .A4(new_n911_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n338_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1352gat));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n920_), .B2(new_n666_), .ZN(new_n927_));
  AOI211_X1 g726(.A(KEYINPUT126), .B(new_n294_), .C1(new_n918_), .C2(new_n919_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n927_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n929_), .ZN(new_n931_));
  AOI21_X1  g730(.A(KEYINPUT123), .B1(new_n893_), .B2(new_n911_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n911_), .ZN(new_n933_));
  NOR4_X1   g732(.A1(new_n824_), .A2(new_n917_), .A3(new_n635_), .A4(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n666_), .B1(new_n932_), .B2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT126), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n920_), .A2(new_n926_), .A3(new_n666_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n931_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n930_), .A2(new_n938_), .ZN(G1353gat));
  OR2_X1    g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  NAND2_X1  g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  AND4_X1   g740(.A1(new_n351_), .A2(new_n920_), .A3(new_n940_), .A4(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n920_), .B2(new_n351_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1354gat));
  AOI21_X1  g743(.A(G218gat), .B1(new_n920_), .B2(new_n627_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n672_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(G218gat), .B2(new_n946_), .ZN(G1355gat));
endmodule


