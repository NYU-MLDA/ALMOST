//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n941_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n969_, new_n970_, new_n971_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n985_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT10), .B(G99gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(G106gat), .ZN(new_n209_));
  AND2_X1   g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  OAI22_X1  g011(.A1(new_n210_), .A2(new_n211_), .B1(KEYINPUT9), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(new_n212_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n213_), .A2(new_n218_), .A3(KEYINPUT64), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT64), .B1(new_n213_), .B2(new_n218_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n207_), .B(new_n209_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n221_));
  OR3_X1    g020(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n205_), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n222_), .B(new_n223_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT66), .B1(new_n210_), .B2(new_n211_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n215_), .A2(new_n228_), .A3(new_n217_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n226_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT8), .ZN(new_n233_));
  INV_X1    g032(.A(new_n223_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT65), .B1(new_n236_), .B2(new_n207_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT8), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n230_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n233_), .A2(KEYINPUT69), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT69), .B1(new_n233_), .B2(new_n239_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n221_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243_));
  INV_X1    g042(.A(G64gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G57gat), .ZN(new_n245_));
  INV_X1    g044(.A(G57gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G64gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G71gat), .B(G78gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n243_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT11), .B1(new_n245_), .B2(new_n247_), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n254_), .A2(KEYINPUT67), .A3(new_n251_), .ZN(new_n255_));
  OAI22_X1  g054(.A1(new_n253_), .A2(new_n255_), .B1(new_n249_), .B2(new_n248_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n243_), .A3(new_n252_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT67), .B1(new_n254_), .B2(new_n251_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n248_), .A2(new_n249_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n261_), .A2(KEYINPUT12), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n242_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n238_), .B1(new_n237_), .B2(new_n230_), .ZN(new_n264_));
  AND4_X1   g063(.A1(new_n231_), .A2(new_n226_), .A3(new_n230_), .A4(new_n238_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n221_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT12), .B1(new_n266_), .B2(new_n261_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n261_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G230gat), .A2(G233gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n263_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n207_), .B1(new_n208_), .B2(G106gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n213_), .A2(new_n218_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n213_), .A2(new_n218_), .A3(KEYINPUT64), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(new_n233_), .B2(new_n239_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n279_), .A2(KEYINPUT68), .A3(new_n260_), .A4(new_n256_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n268_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n266_), .A2(new_n261_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n272_), .B(new_n280_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n271_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G120gat), .B(G148gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT5), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G176gat), .B(G204gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n271_), .A2(new_n284_), .A3(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(KEYINPUT70), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT70), .B1(new_n290_), .B2(new_n292_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n202_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n295_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(KEYINPUT13), .A3(new_n293_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT71), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G232gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT34), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(KEYINPUT35), .ZN(new_n310_));
  INV_X1    g109(.A(G36gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(G29gat), .ZN(new_n312_));
  INV_X1    g111(.A(G29gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(G36gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G50gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(G43gat), .ZN(new_n317_));
  INV_X1    g116(.A(G43gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G50gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n312_), .A2(new_n314_), .A3(new_n317_), .A4(new_n319_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n310_), .B1(new_n279_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT69), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n233_), .A2(new_n239_), .A3(KEYINPUT69), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n278_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n323_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n321_), .A2(new_n322_), .A3(new_n329_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n324_), .B1(new_n328_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n309_), .A2(KEYINPUT35), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n336_), .B(KEYINPUT72), .Z(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n324_), .B(new_n337_), .C1(new_n328_), .C2(new_n334_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT76), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G190gat), .B(G218gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G134gat), .B(G162gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT36), .Z(new_n346_));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n339_), .A2(new_n347_), .A3(new_n340_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n342_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n345_), .A2(KEYINPUT36), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n339_), .A2(new_n350_), .A3(new_n340_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT74), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n339_), .A2(new_n353_), .A3(new_n350_), .A4(new_n340_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n349_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n341_), .A2(new_n346_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT75), .B1(new_n360_), .B2(KEYINPUT37), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n352_), .A2(new_n354_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT37), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n358_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G1gat), .A2(G8gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT14), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G15gat), .A2(G22gat), .ZN(new_n369_));
  AND2_X1   g168(.A1(G15gat), .A2(G22gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(G1gat), .A2(G8gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n367_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G15gat), .B(G22gat), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n375_), .A2(new_n367_), .A3(new_n372_), .A4(new_n368_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G231gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(new_n261_), .ZN(new_n380_));
  XOR2_X1   g179(.A(G127gat), .B(G155gat), .Z(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G183gat), .B(G211gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT17), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n380_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n385_), .A2(new_n386_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n380_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT79), .B1(new_n388_), .B2(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n366_), .A2(new_n396_), .ZN(new_n397_));
  OR3_X1    g196(.A1(new_n307_), .A2(KEYINPUT80), .A3(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT80), .B1(new_n307_), .B2(new_n397_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n407_));
  INV_X1    g206(.A(G141gat), .ZN(new_n408_));
  INV_X1    g207(.A(G148gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT87), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(KEYINPUT87), .A3(new_n407_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n406_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT88), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n403_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n400_), .B1(KEYINPUT1), .B2(new_n402_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(KEYINPUT1), .B2(new_n402_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G141gat), .B(G148gat), .Z(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT29), .B1(new_n419_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G197gat), .B(G204gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT21), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G218gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(G211gat), .ZN(new_n430_));
  INV_X1    g229(.A(G211gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G218gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n427_), .B2(new_n426_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT94), .ZN(new_n436_));
  INV_X1    g235(.A(G197gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(G204gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(G204gat), .ZN(new_n439_));
  INV_X1    g238(.A(G204gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(G197gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(KEYINPUT21), .B(new_n438_), .C1(new_n442_), .C2(new_n436_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT95), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n435_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n435_), .B2(new_n443_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n434_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n425_), .A2(new_n447_), .A3(KEYINPUT93), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G228gat), .A2(G233gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n449_), .B(KEYINPUT92), .Z(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n425_), .A2(new_n447_), .A3(KEYINPUT93), .A4(new_n450_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G78gat), .B(G106gat), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n406_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n402_), .B(new_n401_), .C1(new_n460_), .C2(new_n417_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(new_n423_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT89), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n461_), .A2(new_n465_), .A3(new_n462_), .A4(new_n423_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G22gat), .B(G50gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(KEYINPUT91), .Z(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n459_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT96), .ZN(new_n474_));
  INV_X1    g273(.A(new_n471_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n458_), .A3(new_n469_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n457_), .A2(new_n472_), .A3(new_n474_), .A4(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n472_), .A3(new_n476_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n456_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n473_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G226gat), .A2(G233gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n483_), .B(KEYINPUT19), .Z(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT97), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n435_), .A2(new_n443_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT95), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n435_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n487_), .A2(new_n488_), .B1(new_n433_), .B2(new_n428_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT25), .B(G183gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT26), .B(G190gat), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT24), .ZN(new_n493_));
  INV_X1    g292(.A(G169gat), .ZN(new_n494_));
  INV_X1    g293(.A(G176gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G183gat), .A2(G190gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT23), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(G169gat), .B2(G176gat), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n492_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G183gat), .ZN(new_n505_));
  INV_X1    g304(.A(G190gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n499_), .A2(new_n500_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT99), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n509_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G169gat), .A2(G176gat), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT83), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT98), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(KEYINPUT98), .A3(new_n516_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n494_), .A2(KEYINPUT22), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n494_), .A2(KEYINPUT22), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(G176gat), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n519_), .A2(new_n520_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n504_), .B1(new_n512_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT20), .B1(new_n489_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT84), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n517_), .A2(new_n502_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(new_n492_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n490_), .A2(new_n491_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n530_), .B(KEYINPUT84), .C1(new_n517_), .C2(new_n502_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n501_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n521_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n534_), .A2(KEYINPUT85), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(KEYINPUT85), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n523_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n537_), .A2(new_n515_), .A3(new_n516_), .A4(new_n508_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n533_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(new_n447_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n485_), .B1(new_n526_), .B2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G8gat), .B(G36gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT18), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G64gat), .B(G92gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT20), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n489_), .B2(new_n525_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n539_), .A2(new_n447_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n484_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n541_), .A2(new_n545_), .A3(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n550_), .A2(KEYINPUT27), .ZN(new_n551_));
  INV_X1    g350(.A(new_n545_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n526_), .A2(new_n540_), .A3(new_n485_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n484_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n552_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n524_), .A2(new_n511_), .A3(new_n510_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n504_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT20), .B1(new_n447_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n487_), .A2(new_n488_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n560_), .A2(new_n434_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n484_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n559_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n485_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n546_), .B1(new_n447_), .B2(new_n558_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n560_), .A2(new_n434_), .A3(new_n538_), .A4(new_n533_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n552_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n550_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT27), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n551_), .A2(new_n555_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G1gat), .B(G29gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(G85gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT0), .B(G57gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G127gat), .B(G134gat), .Z(new_n577_));
  XOR2_X1   g376(.A(G113gat), .B(G120gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n461_), .A2(new_n423_), .A3(new_n579_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT4), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT4), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n584_), .B(new_n580_), .C1(new_n419_), .C2(new_n424_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G225gat), .A2(G233gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT100), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n576_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n588_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n594_), .A2(new_n575_), .A3(new_n590_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n482_), .A2(new_n571_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n545_), .A2(KEYINPUT32), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n541_), .A2(new_n598_), .A3(new_n549_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n596_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n581_), .A2(new_n588_), .A3(new_n582_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n576_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT102), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n583_), .A2(new_n593_), .A3(new_n585_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n604_), .A2(new_n576_), .A3(KEYINPUT102), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT33), .B(new_n575_), .C1(new_n594_), .C2(new_n590_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n568_), .A2(new_n610_), .A3(new_n611_), .A4(new_n550_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n575_), .B1(new_n594_), .B2(new_n590_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT101), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(KEYINPUT101), .A3(new_n614_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n603_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n597_), .B1(new_n618_), .B2(new_n482_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G227gat), .A2(G233gat), .ZN(new_n620_));
  INV_X1    g419(.A(G15gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT30), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n539_), .B(new_n624_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n580_), .A2(KEYINPUT31), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n580_), .A2(KEYINPUT31), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(KEYINPUT86), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n539_), .B(new_n623_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n628_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G71gat), .B(G99gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(G43gat), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n630_), .A2(new_n632_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n569_), .A2(new_n570_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n555_), .A2(KEYINPUT27), .A3(new_n550_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n477_), .A2(new_n481_), .A3(new_n638_), .A4(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n635_), .A2(new_n636_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n596_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT103), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n477_), .A2(new_n481_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n596_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n637_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n644_), .A2(new_n646_), .A3(new_n647_), .A4(new_n571_), .ZN(new_n648_));
  AOI22_X1  g447(.A1(new_n619_), .A2(new_n637_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n377_), .A2(KEYINPUT81), .A3(new_n323_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n323_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT81), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n374_), .A2(new_n376_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n650_), .A2(new_n653_), .B1(new_n333_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT82), .ZN(new_n656_));
  NAND2_X1  g455(.A1(G229gat), .A2(G233gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n332_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n329_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n654_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT81), .B1(new_n377_), .B2(new_n323_), .ZN(new_n662_));
  AND4_X1   g461(.A1(KEYINPUT81), .A2(new_n323_), .A3(new_n374_), .A4(new_n376_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n661_), .B(new_n657_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT82), .ZN(new_n665_));
  OAI22_X1  g464(.A1(new_n662_), .A2(new_n663_), .B1(new_n377_), .B2(new_n323_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n657_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n658_), .A2(new_n665_), .A3(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(G169gat), .B(G197gat), .Z(new_n670_));
  XNOR2_X1  g469(.A(G113gat), .B(G141gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n669_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n658_), .A2(new_n665_), .A3(new_n668_), .A4(new_n672_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n649_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n398_), .A2(new_n399_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT38), .ZN(new_n680_));
  INV_X1    g479(.A(G1gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n645_), .A2(new_n681_), .ZN(new_n682_));
  OR3_X1    g481(.A1(new_n679_), .A2(new_n680_), .A3(new_n682_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n302_), .A2(new_n395_), .A3(new_n677_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n649_), .A2(new_n356_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G1gat), .B1(new_n686_), .B2(new_n596_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n680_), .B1(new_n679_), .B2(new_n682_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(new_n687_), .A3(new_n688_), .ZN(G1324gat));
  NOR2_X1   g488(.A1(new_n571_), .A2(G8gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n692_));
  INV_X1    g491(.A(new_n571_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n693_), .A3(new_n685_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n694_), .B2(G8gat), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(G8gat), .A3(new_n692_), .ZN(new_n696_));
  OAI22_X1  g495(.A1(new_n679_), .A2(new_n691_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1325gat));
  OAI21_X1  g498(.A(G15gat), .B1(new_n686_), .B2(new_n637_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT41), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT41), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n641_), .A2(new_n621_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n703_), .B(new_n704_), .C1(new_n679_), .C2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n701_), .B(new_n702_), .C1(new_n679_), .C2(new_n705_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT105), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1326gat));
  XNOR2_X1  g508(.A(new_n644_), .B(KEYINPUT106), .ZN(new_n710_));
  OAI21_X1  g509(.A(G22gat), .B1(new_n686_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT42), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n710_), .A2(G22gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n679_), .B2(new_n713_), .ZN(G1327gat));
  NAND3_X1  g513(.A1(new_n301_), .A2(new_n395_), .A3(new_n676_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n619_), .A2(new_n637_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n643_), .A2(new_n648_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n360_), .A2(KEYINPUT75), .A3(KEYINPUT37), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n363_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n721_), .A2(new_n722_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n717_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n649_), .A2(KEYINPUT43), .A3(new_n366_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n716_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n649_), .B2(new_n366_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n643_), .A2(new_n648_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n617_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n612_), .A2(new_n732_), .A3(new_n615_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n644_), .B1(new_n733_), .B2(new_n603_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n641_), .B1(new_n734_), .B2(new_n597_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n717_), .B(new_n723_), .C1(new_n731_), .C2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n715_), .B1(new_n730_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT107), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n728_), .A2(new_n729_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(KEYINPUT44), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(G29gat), .A3(new_n645_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n356_), .A2(new_n395_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n302_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n678_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n313_), .B1(new_n745_), .B2(new_n596_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n742_), .A2(new_n746_), .ZN(G1328gat));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n739_), .A2(new_n693_), .A3(new_n740_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n311_), .A2(KEYINPUT108), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n571_), .A2(G36gat), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT45), .B1(new_n745_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n744_), .A2(new_n678_), .A3(new_n756_), .A4(new_n752_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n754_), .A2(new_n755_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n748_), .B1(new_n751_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n758_), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT46), .B(new_n760_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1329gat));
  OAI21_X1  g561(.A(new_n318_), .B1(new_n745_), .B2(new_n637_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n641_), .A2(G43gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n737_), .B2(KEYINPUT44), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n739_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n729_), .B1(new_n737_), .B2(KEYINPUT107), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n727_), .B(new_n715_), .C1(new_n730_), .C2(new_n736_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n764_), .B(new_n766_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n763_), .B1(new_n767_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT47), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n763_), .C1(new_n767_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1330gat));
  NAND3_X1  g575(.A1(new_n741_), .A2(G50gat), .A3(new_n482_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n316_), .B1(new_n745_), .B2(new_n710_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1331gat));
  NOR2_X1   g578(.A1(new_n649_), .A2(new_n676_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n781_), .A2(new_n397_), .A3(new_n301_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n246_), .A3(new_n645_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n395_), .A2(new_n676_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n307_), .A2(new_n685_), .A3(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n645_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n786_), .B2(new_n246_), .ZN(G1332gat));
  NOR2_X1   g586(.A1(new_n571_), .A2(G64gat), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT110), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n782_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT48), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n785_), .A2(new_n693_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G64gat), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT48), .B(new_n244_), .C1(new_n785_), .C2(new_n693_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(G1333gat));
  INV_X1    g594(.A(G71gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n782_), .A2(new_n796_), .A3(new_n641_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n785_), .A2(new_n641_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(G71gat), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT49), .B(new_n796_), .C1(new_n785_), .C2(new_n641_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(G1334gat));
  INV_X1    g601(.A(G78gat), .ZN(new_n803_));
  INV_X1    g602(.A(new_n710_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n782_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n785_), .A2(new_n804_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(G78gat), .ZN(new_n808_));
  AOI211_X1 g607(.A(KEYINPUT50), .B(new_n803_), .C1(new_n785_), .C2(new_n804_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n805_), .B1(new_n808_), .B2(new_n809_), .ZN(G1335gat));
  NOR3_X1   g609(.A1(new_n301_), .A2(new_n396_), .A3(new_n676_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n812_), .A2(KEYINPUT112), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(KEYINPUT112), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(G85gat), .B1(new_n815_), .B2(new_n596_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n743_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n307_), .A2(KEYINPUT111), .A3(new_n817_), .A4(new_n780_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n303_), .A2(new_n305_), .A3(new_n817_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n781_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n214_), .A3(new_n645_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n816_), .A2(new_n823_), .ZN(G1336gat));
  OAI21_X1  g623(.A(G92gat), .B1(new_n815_), .B2(new_n571_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n822_), .A2(new_n212_), .A3(new_n693_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1337gat));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(KEYINPUT114), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n637_), .A2(new_n208_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n822_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n637_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n832_));
  INV_X1    g631(.A(G99gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT114), .B1(new_n835_), .B2(new_n828_), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT115), .Z(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n831_), .B(new_n837_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1338gat));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n812_), .A2(new_n644_), .ZN(new_n843_));
  INV_X1    g642(.A(G106gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT116), .B(G106gat), .C1(new_n812_), .C2(new_n644_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(KEYINPUT52), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n842_), .B(new_n848_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n822_), .A2(new_n844_), .A3(new_n482_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT53), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n847_), .A2(new_n853_), .A3(new_n849_), .A4(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1339gat));
  NOR3_X1   g654(.A1(new_n640_), .A2(new_n596_), .A3(new_n637_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n672_), .B1(new_n666_), .B2(new_n657_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n667_), .B1(new_n655_), .B2(KEYINPUT118), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n650_), .A2(new_n653_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n860_), .A2(KEYINPUT118), .A3(new_n661_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n862_), .A2(new_n675_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n292_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT119), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n292_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n270_), .B1(new_n263_), .B2(new_n269_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n271_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n263_), .A2(new_n269_), .A3(KEYINPUT55), .A4(new_n270_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT56), .B1(new_n873_), .B2(new_n289_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n875_));
  AOI211_X1 g674(.A(new_n875_), .B(new_n291_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n868_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n868_), .B(KEYINPUT58), .C1(new_n874_), .C2(new_n876_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n676_), .A2(new_n292_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n863_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n356_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  OAI22_X1  g684(.A1(new_n881_), .A2(new_n366_), .B1(new_n885_), .B2(KEYINPUT57), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(KEYINPUT57), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n395_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n296_), .A2(new_n299_), .A3(new_n784_), .A4(new_n890_), .ZN(new_n891_));
  OR2_X1    g690(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n892_));
  OR3_X1    g691(.A1(new_n723_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  OAI22_X1  g692(.A1(new_n723_), .A2(new_n891_), .B1(KEYINPUT117), .B2(KEYINPUT54), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n857_), .B1(new_n889_), .B2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G113gat), .B1(new_n896_), .B2(new_n676_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT120), .B1(new_n896_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n885_), .A2(KEYINPUT57), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n723_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n887_), .A3(new_n902_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n903_), .A2(new_n395_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n900_), .B(KEYINPUT59), .C1(new_n904_), .C2(new_n857_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n899_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n889_), .A2(new_n895_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(new_n898_), .A3(new_n856_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n676_), .A2(G113gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT121), .Z(new_n911_));
  AOI21_X1  g710(.A(new_n897_), .B1(new_n909_), .B2(new_n911_), .ZN(G1340gat));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913_));
  INV_X1    g712(.A(G120gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n306_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n906_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n896_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT122), .B1(new_n914_), .B2(KEYINPUT60), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n914_), .B1(new_n301_), .B2(KEYINPUT60), .ZN(new_n919_));
  MUX2_X1   g718(.A(KEYINPUT122), .B(new_n918_), .S(new_n919_), .Z(new_n920_));
  NOR2_X1   g719(.A1(new_n917_), .A2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n913_), .B1(new_n916_), .B2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n921_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n908_), .A2(new_n307_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n899_), .B2(new_n905_), .ZN(new_n925_));
  OAI211_X1 g724(.A(KEYINPUT123), .B(new_n923_), .C1(new_n925_), .C2(new_n914_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n922_), .A2(new_n926_), .ZN(G1341gat));
  AOI21_X1  g726(.A(G127gat), .B1(new_n896_), .B2(new_n396_), .ZN(new_n928_));
  INV_X1    g727(.A(G127gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(new_n396_), .B2(KEYINPUT124), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(KEYINPUT124), .B2(new_n929_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n928_), .B1(new_n909_), .B2(new_n931_), .ZN(G1342gat));
  INV_X1    g731(.A(G134gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n896_), .A2(new_n933_), .A3(new_n356_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n906_), .A2(new_n723_), .A3(new_n908_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(new_n933_), .ZN(G1343gat));
  NAND3_X1  g735(.A1(new_n571_), .A2(new_n645_), .A3(new_n637_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n904_), .A2(new_n644_), .A3(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n676_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n307_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n396_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(KEYINPUT61), .B(G155gat), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n943_), .B(new_n944_), .ZN(G1346gat));
  INV_X1    g744(.A(G162gat), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n938_), .A2(new_n946_), .A3(new_n356_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n938_), .A2(new_n723_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n946_), .ZN(G1347gat));
  NAND2_X1  g748(.A1(new_n693_), .A2(new_n646_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n904_), .A2(new_n804_), .A3(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(new_n676_), .ZN(new_n952_));
  OR3_X1    g751(.A1(new_n952_), .A2(new_n534_), .A3(new_n522_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(G169gat), .ZN(new_n954_));
  AND2_X1   g753(.A1(new_n954_), .A2(KEYINPUT62), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n954_), .A2(KEYINPUT62), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n953_), .B1(new_n955_), .B2(new_n956_), .ZN(G1348gat));
  NAND3_X1  g756(.A1(new_n951_), .A2(new_n495_), .A3(new_n302_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n950_), .A2(new_n482_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n907_), .A2(new_n959_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G176gat), .B1(new_n960_), .B2(new_n306_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n958_), .A2(new_n961_), .ZN(G1349gat));
  NOR2_X1   g761(.A1(new_n395_), .A2(new_n490_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n907_), .A2(new_n396_), .A3(new_n959_), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n951_), .A2(new_n963_), .B1(new_n964_), .B2(new_n505_), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n951_), .A2(new_n356_), .A3(new_n491_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n951_), .A2(new_n723_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n966_), .B1(new_n967_), .B2(new_n506_), .ZN(G1351gat));
  NAND4_X1  g767(.A1(new_n693_), .A2(new_n482_), .A3(new_n596_), .A4(new_n637_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n904_), .A2(new_n969_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n970_), .A2(new_n676_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g771(.A1(new_n970_), .A2(new_n307_), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g773(.A(new_n395_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n970_), .A2(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977_));
  NOR2_X1   g776(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(KEYINPUT125), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n976_), .B1(new_n977_), .B2(new_n979_), .ZN(new_n980_));
  XOR2_X1   g779(.A(new_n979_), .B(KEYINPUT126), .Z(new_n981_));
  AOI21_X1  g780(.A(new_n980_), .B1(new_n976_), .B2(new_n981_), .ZN(G1354gat));
  NAND2_X1  g781(.A1(new_n970_), .A2(new_n356_), .ZN(new_n983_));
  XOR2_X1   g782(.A(KEYINPUT127), .B(G218gat), .Z(new_n984_));
  NOR2_X1   g783(.A1(new_n366_), .A2(new_n984_), .ZN(new_n985_));
  AOI22_X1  g784(.A1(new_n983_), .A2(new_n984_), .B1(new_n970_), .B2(new_n985_), .ZN(G1355gat));
endmodule


