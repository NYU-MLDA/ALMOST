//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_, new_n976_;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT78), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT78), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G169gat), .A3(G176gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT25), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT25), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT26), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT26), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G190gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n212_), .A2(new_n214_), .A3(new_n216_), .A4(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT23), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n210_), .A2(new_n219_), .A3(new_n224_), .A4(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n220_), .A2(new_n222_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n211_), .A2(new_n215_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G169gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT22), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT22), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n232_), .A2(new_n238_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n228_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G211gat), .B(G218gat), .Z(new_n241_));
  NOR2_X1   g040(.A1(G197gat), .A2(G204gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G197gat), .A2(G204gat), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n241_), .A2(KEYINPUT21), .A3(new_n243_), .A4(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(KEYINPUT21), .A3(new_n244_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT21), .ZN(new_n247_));
  AND2_X1   g046(.A1(G197gat), .A2(G204gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(new_n242_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G211gat), .B(G218gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT20), .B1(new_n240_), .B2(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n208_), .B1(G169gat), .B2(G176gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n206_), .A2(KEYINPUT78), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT86), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT86), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n207_), .A2(new_n209_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n254_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT87), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n232_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT87), .B1(G183gat), .B2(G190gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n224_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n260_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n233_), .A2(new_n237_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT24), .A3(new_n206_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n219_), .A2(new_n224_), .A3(new_n227_), .A4(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n205_), .A2(new_n206_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n273_), .A2(KEYINPUT85), .A3(new_n219_), .A4(new_n227_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n267_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n253_), .B1(new_n252_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G226gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT19), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n245_), .A2(new_n251_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n267_), .A2(new_n281_), .A3(new_n270_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT20), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(new_n240_), .B2(new_n252_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n278_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT91), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n203_), .B1(new_n287_), .B2(new_n294_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n267_), .A2(new_n281_), .A3(new_n272_), .A4(new_n274_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n279_), .A3(new_n284_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT89), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n296_), .A2(KEYINPUT89), .A3(new_n284_), .A4(new_n279_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n272_), .A2(new_n274_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n207_), .A2(new_n209_), .A3(new_n258_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n258_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n238_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n261_), .A2(new_n232_), .B1(new_n224_), .B2(new_n264_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n252_), .B1(new_n303_), .B2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n228_), .A2(new_n239_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n283_), .B1(new_n310_), .B2(new_n281_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n302_), .B1(new_n312_), .B2(new_n278_), .ZN(new_n313_));
  AOI211_X1 g112(.A(KEYINPUT88), .B(new_n279_), .C1(new_n309_), .C2(new_n311_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n301_), .B(new_n293_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n295_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT92), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n301_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n294_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT88), .B1(new_n276_), .B2(new_n279_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n312_), .A2(new_n302_), .A3(new_n278_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n324_), .A2(KEYINPUT92), .A3(new_n293_), .A4(new_n301_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n319_), .A2(new_n321_), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n317_), .B1(new_n326_), .B2(new_n203_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT81), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT3), .ZN(new_n331_));
  NOR3_X1   g130(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n331_), .A2(new_n334_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G155gat), .ZN(new_n340_));
  INV_X1    g139(.A(G162gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(KEYINPUT80), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(G155gat), .B2(G162gat), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n342_), .A2(new_n344_), .B1(G155gat), .B2(G162gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n344_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT1), .B1(new_n340_), .B2(new_n341_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(G155gat), .A3(G162gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G141gat), .B(G148gat), .Z(new_n351_));
  AOI22_X1  g150(.A1(new_n339_), .A2(new_n345_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G127gat), .B(G134gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G113gat), .B(G120gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n356_), .A3(KEYINPUT93), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n337_), .B(new_n338_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n330_), .A2(KEYINPUT3), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n345_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n342_), .A2(new_n344_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n347_), .A2(new_n349_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n351_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n363_), .A3(KEYINPUT93), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n355_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n357_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n357_), .B2(new_n365_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n360_), .A2(new_n363_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(new_n356_), .A3(new_n369_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n367_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n368_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G57gat), .B(G85gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n368_), .B(new_n380_), .C1(new_n370_), .C2(new_n374_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G22gat), .B(G50gat), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n360_), .A2(new_n363_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT28), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT28), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n360_), .A2(new_n363_), .A3(new_n391_), .A4(new_n387_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n389_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n386_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(new_n352_), .B2(new_n387_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n392_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT82), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n389_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n385_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(new_n400_), .A3(KEYINPUT84), .ZN(new_n401_));
  XOR2_X1   g200(.A(G78gat), .B(G106gat), .Z(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n395_), .A2(new_n400_), .A3(KEYINPUT84), .A4(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n395_), .A2(new_n400_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n252_), .B1(new_n352_), .B2(new_n387_), .ZN(new_n410_));
  AND2_X1   g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n410_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n409_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n406_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n416_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(new_n405_), .A3(new_n403_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n384_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n287_), .A2(new_n293_), .A3(KEYINPUT32), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n293_), .A2(KEYINPUT32), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n384_), .B(new_n423_), .C1(new_n320_), .C2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n370_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n372_), .A2(new_n367_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT96), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT96), .B1(new_n370_), .B2(new_n427_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n380_), .B1(new_n366_), .B2(new_n373_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT95), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n383_), .A2(new_n435_), .A3(KEYINPUT33), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT33), .B1(new_n383_), .B2(new_n435_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n434_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n425_), .B1(new_n326_), .B2(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n420_), .A2(new_n405_), .A3(new_n403_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n403_), .A2(new_n405_), .B1(new_n409_), .B2(new_n417_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n327_), .A2(new_n422_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445_));
  INV_X1    g244(.A(G15gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT30), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT31), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G71gat), .B(G99gat), .ZN(new_n450_));
  INV_X1    g249(.A(G43gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n240_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n449_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT79), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n455_), .A2(new_n356_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n356_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n202_), .B1(new_n444_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n457_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n422_), .A2(new_n327_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n419_), .A2(new_n421_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n383_), .A2(new_n435_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n465_), .A2(new_n436_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n466_), .A2(new_n319_), .A3(new_n321_), .A4(new_n325_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n462_), .B1(new_n467_), .B2(new_n425_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT97), .B(new_n460_), .C1(new_n461_), .C2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n326_), .A2(new_n203_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n316_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n471_), .A2(new_n462_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n460_), .A2(new_n384_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n459_), .A2(new_n469_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G232gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT34), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT35), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT10), .B(G99gat), .Z(new_n483_));
  INV_X1    g282(.A(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G85gat), .B(G92gat), .Z(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT9), .ZN(new_n487_));
  INV_X1    g286(.A(G85gat), .ZN(new_n488_));
  INV_X1    g287(.A(G92gat), .ZN(new_n489_));
  OR3_X1    g288(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT9), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT6), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n485_), .A2(new_n487_), .A3(new_n490_), .A4(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  OR3_X1    g293(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n492_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n497_), .A2(KEYINPUT64), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n496_), .A2(new_n486_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n498_), .B1(new_n496_), .B2(new_n486_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n493_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G29gat), .B(G36gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT15), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT66), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n501_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n509_), .A2(new_n504_), .B1(new_n480_), .B2(new_n479_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n482_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n506_), .A2(new_n507_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT66), .B1(new_n501_), .B2(new_n505_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n510_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(new_n481_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT69), .B1(new_n511_), .B2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(new_n482_), .A3(new_n510_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n481_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G190gat), .B(G218gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(G134gat), .B(G162gat), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n522_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n523_), .A2(KEYINPUT36), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT36), .B1(new_n523_), .B2(new_n524_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n516_), .A2(new_n520_), .A3(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n526_), .B(KEYINPUT67), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n517_), .A2(new_n518_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n476_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT12), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT65), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n537_));
  XOR2_X1   g336(.A(G71gat), .B(G78gat), .Z(new_n538_));
  OR2_X1    g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n538_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n496_), .A2(new_n486_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n498_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n496_), .A2(new_n486_), .A3(new_n498_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n542_), .B1(new_n547_), .B2(new_n493_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n542_), .B(new_n493_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n535_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n542_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n534_), .A2(KEYINPUT65), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n501_), .A2(new_n553_), .B1(new_n554_), .B2(new_n535_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n552_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n558_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G120gat), .B(G148gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT5), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n557_), .A2(new_n559_), .A3(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n565_), .A2(KEYINPUT13), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT13), .B1(new_n565_), .B2(new_n567_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n542_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT72), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT70), .B(G8gat), .ZN(new_n575_));
  INV_X1    g374(.A(G1gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT14), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G15gat), .B(G22gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT71), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(new_n581_), .A3(new_n578_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G1gat), .B(G8gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n582_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n584_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n574_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT72), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n573_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G127gat), .B(G155gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT17), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n590_), .A2(new_n594_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n599_), .B(KEYINPUT17), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n590_), .B2(new_n594_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n589_), .A2(new_n505_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n585_), .A2(new_n588_), .A3(new_n504_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G229gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT75), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n608_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT76), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT76), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n608_), .A2(new_n614_), .A3(new_n609_), .A4(new_n611_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n609_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n504_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n617_));
  OAI211_X1 g416(.A(G229gat), .B(G233gat), .C1(new_n616_), .C2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n613_), .A2(new_n615_), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G113gat), .B(G141gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G169gat), .B(G197gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n620_), .B(new_n621_), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n613_), .A2(new_n615_), .A3(new_n618_), .A4(new_n622_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n571_), .A2(new_n607_), .A3(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n533_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n384_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G1gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n626_), .B(KEYINPUT77), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT37), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n531_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT74), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n602_), .A2(new_n605_), .A3(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n592_), .A2(new_n593_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n574_), .A2(new_n589_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n603_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n590_), .A2(new_n594_), .A3(new_n601_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT74), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n527_), .B(KEYINPUT68), .Z(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(KEYINPUT37), .A3(new_n530_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n634_), .A2(new_n570_), .A3(new_n642_), .A4(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n475_), .A2(new_n632_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n475_), .A2(KEYINPUT98), .A3(new_n647_), .A4(new_n632_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n384_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(G1gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n651_), .A3(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n655_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n650_), .A2(new_n651_), .A3(new_n653_), .A4(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n631_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT100), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n631_), .A2(new_n659_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1324gat));
  NAND4_X1  g463(.A1(new_n475_), .A2(new_n471_), .A3(new_n531_), .A4(new_n628_), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT102), .B(KEYINPUT39), .C1(new_n665_), .C2(G8gat), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n665_), .A2(G8gat), .ZN(new_n667_));
  XOR2_X1   g466(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n471_), .A2(new_n575_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n650_), .A2(new_n651_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n650_), .A2(KEYINPUT101), .A3(new_n651_), .A4(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n669_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n669_), .A2(new_n675_), .A3(KEYINPUT40), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1325gat));
  NAND2_X1  g479(.A1(new_n629_), .A2(new_n458_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT41), .B1(new_n681_), .B2(G15gat), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n458_), .A2(new_n446_), .ZN(new_n684_));
  OAI22_X1  g483(.A1(new_n682_), .A2(new_n683_), .B1(new_n648_), .B2(new_n684_), .ZN(G1326gat));
  OR3_X1    g484(.A1(new_n648_), .A2(G22gat), .A3(new_n443_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n629_), .A2(new_n462_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G22gat), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT42), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT42), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(G1327gat));
  INV_X1    g490(.A(KEYINPUT77), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n626_), .B(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n476_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n635_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n639_), .A2(KEYINPUT74), .A3(new_n640_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n532_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n571_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n694_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G29gat), .B1(new_n700_), .B2(new_n384_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n571_), .A2(new_n642_), .A3(new_n627_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n634_), .A2(new_n645_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n475_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n475_), .B2(new_n704_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT44), .B(new_n702_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n707_), .A2(G29gat), .A3(new_n384_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n701_), .B1(new_n708_), .B2(new_n711_), .ZN(G1328gat));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713_));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n702_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n422_), .A2(new_n327_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n440_), .A2(new_n443_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n458_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n474_), .B1(new_n718_), .B2(KEYINPUT97), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n444_), .A2(new_n202_), .A3(new_n458_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n704_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT43), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n475_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n715_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n327_), .B1(new_n724_), .B2(KEYINPUT44), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n714_), .B1(new_n725_), .B2(new_n711_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n694_), .A2(new_n714_), .A3(new_n471_), .A4(new_n699_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT103), .Z(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n727_), .B(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n713_), .B1(new_n726_), .B2(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n724_), .A2(KEYINPUT44), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n707_), .A2(new_n471_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G36gat), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n727_), .B(new_n729_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(KEYINPUT46), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n732_), .A2(new_n737_), .ZN(G1329gat));
  NAND4_X1  g537(.A1(new_n475_), .A2(new_n458_), .A3(new_n632_), .A4(new_n699_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n451_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT105), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n707_), .A2(G43gat), .A3(new_n458_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(new_n733_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT47), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n741_), .B(new_n745_), .C1(new_n742_), .C2(new_n733_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1330gat));
  INV_X1    g546(.A(G50gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n700_), .A2(new_n748_), .A3(new_n462_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n707_), .A2(new_n462_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n733_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G50gat), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n733_), .A2(new_n751_), .A3(new_n750_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n749_), .B1(new_n753_), .B2(new_n754_), .ZN(G1331gat));
  AOI21_X1  g554(.A(KEYINPUT37), .B1(new_n528_), .B2(new_n530_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n645_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n756_), .A2(new_n697_), .A3(new_n757_), .ZN(new_n758_));
  AND4_X1   g557(.A1(new_n475_), .A2(new_n627_), .A3(new_n571_), .A4(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(G57gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n384_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n632_), .A2(new_n570_), .A3(new_n697_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n533_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n533_), .A2(KEYINPUT107), .A3(new_n762_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n384_), .A3(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n761_), .B1(new_n767_), .B2(new_n760_), .ZN(G1332gat));
  INV_X1    g567(.A(G64gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n759_), .A2(new_n769_), .A3(new_n471_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n765_), .A2(new_n471_), .A3(new_n766_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(G64gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G64gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1333gat));
  INV_X1    g574(.A(G71gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n759_), .A2(new_n776_), .A3(new_n458_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n765_), .A2(new_n458_), .A3(new_n766_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(G71gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G71gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1334gat));
  INV_X1    g581(.A(G78gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n759_), .A2(new_n783_), .A3(new_n462_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n765_), .A2(new_n462_), .A3(new_n766_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(G78gat), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n785_), .B2(G78gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(G1335gat));
  NAND3_X1  g588(.A1(new_n571_), .A2(new_n627_), .A3(new_n697_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT109), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(G85gat), .B1(new_n794_), .B2(new_n652_), .ZN(new_n795_));
  NOR4_X1   g594(.A1(new_n476_), .A2(new_n626_), .A3(new_n570_), .A4(new_n698_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n488_), .A3(new_n384_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1336gat));
  OAI21_X1  g597(.A(G92gat), .B1(new_n794_), .B2(new_n327_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n489_), .A3(new_n471_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n792_), .B2(new_n460_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n796_), .A2(new_n458_), .A3(new_n483_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g604(.A1(new_n796_), .A2(new_n484_), .A3(new_n462_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n462_), .B(new_n791_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n807_), .A2(new_n808_), .A3(G106gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n807_), .B2(G106gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT53), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(new_n806_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1339gat));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n646_), .B2(new_n632_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n758_), .A2(new_n817_), .A3(new_n570_), .A4(new_n693_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT113), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n551_), .A2(KEYINPUT55), .A3(new_n552_), .A4(new_n556_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n501_), .A2(new_n553_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n823_), .A2(new_n549_), .B1(KEYINPUT65), .B2(new_n534_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n558_), .B1(new_n824_), .B2(new_n555_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n824_), .A2(new_n558_), .A3(new_n555_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n829_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n557_), .A2(KEYINPUT112), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n826_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n821_), .B1(new_n833_), .B2(new_n566_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n826_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n557_), .A2(KEYINPUT112), .A3(new_n831_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT112), .B1(new_n557_), .B2(new_n831_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n821_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n564_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n567_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n834_), .A2(new_n840_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n565_), .A2(new_n567_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n611_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n608_), .A2(new_n609_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n846_), .B(new_n623_), .C1(new_n847_), .C2(new_n611_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n625_), .A2(new_n845_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n845_), .B1(new_n625_), .B2(new_n848_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n844_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n843_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n531_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n532_), .B1(new_n843_), .B2(new_n851_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT115), .B1(new_n857_), .B2(KEYINPUT57), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(KEYINPUT57), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT56), .B1(new_n833_), .B2(new_n566_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n838_), .A2(new_n820_), .A3(new_n564_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n567_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n860_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n625_), .A2(new_n848_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT114), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n625_), .A2(new_n845_), .A3(new_n848_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n841_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n869_), .A2(KEYINPUT58), .A3(new_n861_), .A4(new_n862_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n865_), .A2(new_n870_), .A3(new_n704_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n856_), .A2(new_n858_), .A3(new_n859_), .A4(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n819_), .B1(new_n872_), .B2(new_n607_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n472_), .A2(new_n384_), .A3(new_n458_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT116), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT59), .B1(new_n873_), .B2(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n871_), .A2(new_n859_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n853_), .A2(new_n855_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n642_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n875_), .B(new_n878_), .C1(new_n881_), .C2(new_n819_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT118), .B(G113gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n693_), .A2(new_n883_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n877_), .A2(new_n882_), .A3(new_n884_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n873_), .A2(new_n627_), .A3(new_n876_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(G113gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT119), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n877_), .A2(new_n882_), .A3(new_n884_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n889_), .B(new_n890_), .C1(G113gat), .C2(new_n886_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n891_), .ZN(G1340gat));
  NAND2_X1  g691(.A1(new_n877_), .A2(new_n882_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G120gat), .B1(new_n893_), .B2(new_n570_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n873_), .A2(new_n876_), .ZN(new_n895_));
  INV_X1    g694(.A(G120gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n570_), .B2(KEYINPUT60), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n895_), .B(new_n897_), .C1(KEYINPUT60), .C2(new_n896_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n898_), .ZN(G1341gat));
  AOI21_X1  g698(.A(G127gat), .B1(new_n895_), .B2(new_n642_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n893_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT120), .B(G127gat), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n607_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(G1342gat));
  AOI21_X1  g703(.A(G134gat), .B1(new_n895_), .B2(new_n532_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n704_), .A2(G134gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT121), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n901_), .B2(new_n907_), .ZN(G1343gat));
  NAND2_X1  g707(.A1(new_n872_), .A2(new_n607_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n819_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n458_), .A2(new_n471_), .A3(new_n652_), .A4(new_n443_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n626_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g715(.A1(new_n913_), .A2(new_n570_), .ZN(new_n917_));
  XOR2_X1   g716(.A(KEYINPUT122), .B(G148gat), .Z(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1345gat));
  NAND2_X1  g718(.A1(new_n914_), .A2(new_n642_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT61), .B(G155gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1346gat));
  NOR2_X1   g721(.A1(new_n756_), .A2(new_n757_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G162gat), .B1(new_n913_), .B2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n532_), .A2(new_n341_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n913_), .B2(new_n925_), .ZN(G1347gat));
  AOI21_X1  g725(.A(new_n233_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n881_), .A2(new_n819_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n473_), .A2(new_n471_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(new_n627_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT123), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n443_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n927_), .B1(new_n928_), .B2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n934_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n929_), .A2(new_n462_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n937_), .B1(new_n881_), .B2(new_n819_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n626_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n935_), .B(new_n936_), .C1(new_n938_), .C2(new_n939_), .ZN(G1348gat));
  OAI21_X1  g739(.A(new_n237_), .B1(new_n938_), .B2(new_n570_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n911_), .A2(new_n443_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n929_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n943_), .A2(G176gat), .A3(new_n571_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n941_), .B1(new_n942_), .B2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(KEYINPUT125), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n941_), .B(new_n947_), .C1(new_n942_), .C2(new_n944_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(G1349gat));
  AOI211_X1 g748(.A(new_n607_), .B(new_n938_), .C1(new_n212_), .C2(new_n214_), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n911_), .A2(new_n443_), .A3(new_n642_), .A4(new_n943_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n951_), .B2(new_n211_), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n938_), .B2(new_n923_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n532_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n954_));
  XOR2_X1   g753(.A(new_n954_), .B(KEYINPUT126), .Z(new_n955_));
  OAI21_X1  g754(.A(new_n953_), .B1(new_n938_), .B2(new_n955_), .ZN(G1351gat));
  AND4_X1   g755(.A1(new_n460_), .A2(new_n911_), .A3(new_n471_), .A4(new_n422_), .ZN(new_n957_));
  AND3_X1   g756(.A1(new_n957_), .A2(G197gat), .A3(new_n626_), .ZN(new_n958_));
  AOI21_X1  g757(.A(G197gat), .B1(new_n957_), .B2(new_n626_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n957_), .A2(new_n571_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(G204gat), .ZN(new_n962_));
  INV_X1    g761(.A(G204gat), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n957_), .A2(new_n963_), .A3(new_n571_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n964_), .ZN(G1353gat));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n966_));
  INV_X1    g765(.A(G211gat), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n606_), .B1(new_n966_), .B2(new_n967_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(KEYINPUT127), .ZN(new_n970_));
  AND3_X1   g769(.A1(new_n957_), .A2(new_n968_), .A3(new_n970_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n968_), .B1(new_n957_), .B2(new_n970_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n971_), .A2(new_n972_), .ZN(G1354gat));
  INV_X1    g772(.A(G218gat), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n957_), .A2(new_n974_), .A3(new_n532_), .ZN(new_n975_));
  AND2_X1   g774(.A1(new_n957_), .A2(new_n704_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n975_), .B1(new_n976_), .B2(new_n974_), .ZN(G1355gat));
endmodule


