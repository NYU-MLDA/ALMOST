//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G1gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT76), .B(G8gat), .ZN(new_n208_));
  OAI211_X1 g007(.A(G1gat), .B(new_n202_), .C1(new_n208_), .C2(new_n203_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n206_), .A2(new_n209_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G8gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n215_), .A2(KEYINPUT15), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(KEYINPUT15), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n210_), .B(new_n212_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n210_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n215_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(KEYINPUT80), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n224_));
  XOR2_X1   g023(.A(G43gat), .B(G50gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(new_n213_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n212_), .A2(new_n210_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n212_), .B2(new_n210_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n224_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(KEYINPUT79), .A3(new_n227_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n221_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n222_), .A2(KEYINPUT80), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n223_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236_));
  INV_X1    g035(.A(G197gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT81), .B(G169gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n240_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n223_), .A2(new_n233_), .A3(new_n234_), .A4(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G57gat), .ZN(new_n245_));
  INV_X1    g044(.A(G64gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G57gat), .A2(G64gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G71gat), .A2(G78gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G71gat), .A2(G78gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n250_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT67), .ZN(new_n255_));
  AND2_X1   g054(.A1(G57gat), .A2(G64gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G57gat), .A2(G64gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(new_n248_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n250_), .A2(new_n260_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n255_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n259_), .B1(new_n255_), .B2(new_n261_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G85gat), .B(G92gat), .Z(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT9), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G99gat), .A2(G106gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G106gat), .ZN(new_n272_));
  INV_X1    g071(.A(G99gat), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n273_), .A2(KEYINPUT10), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(KEYINPUT10), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n272_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G85gat), .ZN(new_n277_));
  INV_X1    g076(.A(G92gat), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n277_), .A2(new_n278_), .A3(KEYINPUT9), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n266_), .A2(new_n271_), .A3(new_n276_), .A4(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n281_));
  AOI211_X1 g080(.A(G99gat), .B(G106gat), .C1(new_n281_), .C2(KEYINPUT65), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT7), .B1(new_n283_), .B2(KEYINPUT66), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n271_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT8), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n285_), .A2(new_n286_), .A3(new_n265_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n285_), .B2(new_n265_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n280_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n264_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n259_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n252_), .B1(new_n258_), .B2(new_n248_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n260_), .B1(new_n292_), .B2(new_n251_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n261_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n291_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n255_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AND4_X1   g096(.A1(new_n266_), .A2(new_n271_), .A3(new_n276_), .A4(new_n279_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n269_), .A2(new_n270_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n283_), .A2(KEYINPUT66), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n281_), .A2(KEYINPUT65), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(new_n273_), .A3(new_n272_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n299_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n265_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT8), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n285_), .A2(new_n286_), .A3(new_n265_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n298_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n297_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n290_), .A2(new_n310_), .A3(KEYINPUT12), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT12), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n264_), .A2(new_n289_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G230gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT64), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n290_), .A2(new_n310_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n316_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G120gat), .B(G148gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(G204gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT5), .B(G176gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n318_), .A2(new_n320_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n329_), .B(KEYINPUT13), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT68), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G1gat), .B(G29gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(new_n277_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT0), .B(G57gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n334_), .B(new_n335_), .Z(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT2), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n339_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT85), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G155gat), .B(G162gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n339_), .A2(KEYINPUT85), .A3(new_n340_), .A4(new_n343_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n348_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n346_), .A2(new_n349_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n341_), .B(KEYINPUT84), .Z(new_n353_));
  OR2_X1    g152(.A1(new_n347_), .A2(KEYINPUT1), .ZN(new_n354_));
  NAND3_X1  g153(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n338_), .A4(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G127gat), .B(G134gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G113gat), .B(G120gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT91), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n352_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(KEYINPUT4), .A4(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n362_), .A2(KEYINPUT4), .A3(new_n364_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT91), .B1(new_n362_), .B2(KEYINPUT4), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n362_), .A2(new_n369_), .A3(new_n364_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n337_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  AOI211_X1 g173(.A(new_n372_), .B(new_n336_), .C1(new_n368_), .C2(new_n370_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT19), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G211gat), .B(G218gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(G197gat), .B(G204gat), .Z(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(KEYINPUT21), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT88), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT89), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n384_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT21), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n384_), .B(KEYINPUT21), .C1(new_n382_), .C2(new_n385_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n388_), .B(new_n389_), .C1(new_n384_), .C2(new_n382_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n383_), .B1(new_n390_), .B2(new_n381_), .ZN(new_n391_));
  INV_X1    g190(.A(G169gat), .ZN(new_n392_));
  INV_X1    g191(.A(G176gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT22), .B(G169gat), .Z(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n396_), .B2(G176gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G183gat), .A2(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT23), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT23), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(G183gat), .A3(G190gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT83), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(KEYINPUT83), .B2(new_n402_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G183gat), .A2(G190gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n398_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G169gat), .A2(G176gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n409_), .B(KEYINPUT82), .Z(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(KEYINPUT24), .A3(new_n395_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n409_), .B(KEYINPUT82), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT24), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT25), .B(G183gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT26), .B(G190gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n411_), .A2(new_n414_), .A3(new_n403_), .A4(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n408_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n391_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n411_), .A2(new_n417_), .A3(new_n414_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n404_), .A2(new_n407_), .ZN(new_n422_));
  OAI22_X1  g221(.A1(new_n421_), .A2(new_n406_), .B1(new_n397_), .B2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n391_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT90), .ZN(new_n425_));
  OAI211_X1 g224(.A(KEYINPUT20), .B(new_n420_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n391_), .A2(new_n423_), .A3(KEYINPUT90), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n380_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n391_), .A2(new_n419_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n391_), .B2(new_n423_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n379_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT32), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G92gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT18), .B(G64gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n436_), .B(new_n437_), .Z(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n433_), .B1(new_n434_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n429_), .A2(new_n380_), .A3(new_n431_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT94), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n420_), .A2(KEYINPUT20), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n379_), .B1(new_n444_), .B2(new_n424_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n429_), .A2(new_n431_), .A3(KEYINPUT94), .A4(new_n380_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(KEYINPUT32), .A3(new_n438_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n377_), .A2(new_n440_), .A3(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n433_), .B(new_n439_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT33), .B1(new_n375_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n368_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT93), .B1(new_n453_), .B2(new_n370_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n362_), .A2(new_n370_), .A3(new_n364_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT93), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n368_), .A2(new_n456_), .A3(new_n369_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n454_), .A2(new_n336_), .A3(new_n455_), .A4(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n371_), .A2(new_n373_), .A3(new_n337_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT92), .A3(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n450_), .A2(new_n452_), .A3(new_n458_), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n449_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n419_), .A2(KEYINPUT30), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n419_), .A2(KEYINPUT30), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n361_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n419_), .A2(KEYINPUT30), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n419_), .A2(KEYINPUT30), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n360_), .A3(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G15gat), .B(G43gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT31), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n470_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n467_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(new_n473_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n475_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n470_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n466_), .A3(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G228gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n485_), .A2(G228gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(G233gat), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n391_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n492_), .B1(new_n352_), .B2(new_n356_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n490_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G22gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n493_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n391_), .A3(new_n489_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G78gat), .B(G106gat), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n494_), .A2(new_n497_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G22gat), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n503_), .B1(new_n505_), .B2(new_n498_), .ZN(new_n506_));
  INV_X1    g305(.A(G50gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n352_), .A2(new_n492_), .A3(new_n356_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n508_), .A2(KEYINPUT28), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(KEYINPUT28), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n507_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n509_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n512_));
  OAI22_X1  g311(.A1(new_n502_), .A2(new_n506_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n501_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n512_), .A2(new_n511_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n505_), .A2(new_n503_), .A3(new_n498_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n463_), .A2(new_n484_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT95), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n447_), .A2(new_n520_), .A3(new_n439_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n433_), .A2(new_n438_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n520_), .B1(new_n447_), .B2(new_n439_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT27), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT27), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n450_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n479_), .A2(new_n483_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n517_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n515_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n484_), .A2(new_n513_), .A3(new_n517_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n528_), .B(new_n376_), .C1(new_n533_), .C2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n519_), .A2(new_n536_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n215_), .B(new_n280_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT34), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(KEYINPUT35), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT70), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(KEYINPUT70), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n538_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n216_), .A2(new_n217_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(new_n309_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n540_), .A2(KEYINPUT35), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n544_), .B(new_n547_), .C1(KEYINPUT69), .C2(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G134gat), .B(G162gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G190gat), .B(G218gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT36), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n538_), .A2(KEYINPUT69), .A3(new_n542_), .A4(new_n543_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n548_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n538_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n557_), .B(new_n558_), .C1(new_n559_), .C2(new_n546_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n549_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n554_), .B(KEYINPUT36), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n549_), .B2(new_n560_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n561_), .B1(new_n564_), .B2(KEYINPUT73), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n549_), .A2(new_n560_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n566_), .A2(KEYINPUT73), .A3(new_n562_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT37), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n549_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(new_n564_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT74), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT74), .ZN(new_n573_));
  NOR4_X1   g372(.A1(new_n569_), .A2(new_n564_), .A3(new_n573_), .A4(KEYINPUT37), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n568_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT75), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n570_), .A2(KEYINPUT74), .A3(new_n571_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n566_), .A2(new_n562_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(new_n571_), .A3(new_n561_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n573_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(KEYINPUT75), .A3(new_n568_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n577_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n219_), .B(new_n585_), .Z(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n588_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n264_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593_));
  INV_X1    g392(.A(G211gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT16), .B(G183gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n589_), .A2(new_n297_), .A3(new_n590_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n592_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n597_), .A2(new_n598_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n592_), .B2(new_n600_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n584_), .A2(new_n604_), .ZN(new_n605_));
  AND4_X1   g404(.A1(new_n244_), .A2(new_n332_), .A3(new_n537_), .A4(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n205_), .A3(new_n377_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n330_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n604_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n244_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n570_), .B1(new_n519_), .B2(new_n536_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n613_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT98), .Z(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(new_n377_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n609_), .B1(new_n619_), .B2(new_n205_), .ZN(G1324gat));
  INV_X1    g419(.A(new_n208_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n528_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n606_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT99), .ZN(new_n624_));
  OAI21_X1  g423(.A(G8gat), .B1(new_n617_), .B2(new_n528_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT39), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g427(.A(G15gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n618_), .B2(new_n529_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT41), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n606_), .A2(new_n629_), .A3(new_n529_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(new_n518_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n495_), .B1(new_n618_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT42), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n606_), .A2(new_n495_), .A3(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1327gat));
  INV_X1    g438(.A(new_n570_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n519_), .B2(new_n536_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n244_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n330_), .A2(new_n611_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(G29gat), .B1(new_n645_), .B2(new_n377_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n537_), .A2(new_n584_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT43), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n537_), .A2(new_n650_), .A3(new_n584_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n647_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n654_), .B1(new_n652_), .B2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n377_), .A2(G29gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n646_), .B1(new_n657_), .B2(new_n658_), .ZN(G1328gat));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n644_), .A2(G36gat), .A3(new_n528_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT45), .Z(new_n662_));
  AOI21_X1  g461(.A(new_n650_), .B1(new_n537_), .B2(new_n584_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n577_), .A2(new_n583_), .ZN(new_n664_));
  AOI211_X1 g463(.A(KEYINPUT43), .B(new_n664_), .C1(new_n519_), .C2(new_n536_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n643_), .B(new_n656_), .C1(new_n663_), .C2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n666_), .B(new_n622_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G36gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n660_), .B1(new_n662_), .B2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT102), .B(KEYINPUT46), .Z(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(G1329gat));
  OAI211_X1 g470(.A(new_n666_), .B(new_n529_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G43gat), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n484_), .A2(G43gat), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n644_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT103), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n673_), .A2(new_n679_), .A3(new_n676_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(KEYINPUT47), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT47), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n679_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT103), .B(new_n675_), .C1(new_n672_), .C2(G43gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n681_), .A2(new_n685_), .ZN(G1330gat));
  NAND3_X1  g485(.A1(new_n645_), .A2(new_n507_), .A3(new_n634_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n666_), .B(new_n634_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(new_n689_), .A3(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n688_), .B2(G50gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1331gat));
  NOR2_X1   g491(.A1(new_n604_), .A2(new_n244_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n615_), .A2(new_n331_), .A3(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT105), .B(G57gat), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n694_), .A2(new_n376_), .A3(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT106), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n664_), .A2(new_n693_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n537_), .A2(new_n698_), .A3(new_n330_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n245_), .B1(new_n699_), .B2(new_n376_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT107), .Z(G1332gat));
  OAI21_X1  g501(.A(G64gat), .B1(new_n694_), .B2(new_n528_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT48), .ZN(new_n704_));
  INV_X1    g503(.A(new_n699_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n246_), .A3(new_n622_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1333gat));
  OR3_X1    g506(.A1(new_n699_), .A2(G71gat), .A3(new_n484_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n615_), .A2(new_n529_), .A3(new_n331_), .A4(new_n693_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(G71gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G71gat), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT49), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n711_), .A2(new_n712_), .A3(KEYINPUT49), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n708_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(G1334gat));
  OAI21_X1  g518(.A(G78gat), .B1(new_n694_), .B2(new_n518_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT50), .Z(new_n721_));
  NOR3_X1   g520(.A1(new_n699_), .A2(G78gat), .A3(new_n518_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1335gat));
  NOR2_X1   g522(.A1(new_n611_), .A2(new_n244_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n641_), .A2(new_n331_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G85gat), .B1(new_n725_), .B2(new_n377_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n649_), .A2(new_n651_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n727_), .A2(new_n330_), .A3(new_n724_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n376_), .A2(new_n277_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(G1336gat));
  AOI21_X1  g529(.A(G92gat), .B1(new_n725_), .B2(new_n622_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n528_), .A2(new_n278_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n728_), .B2(new_n732_), .ZN(G1337gat));
  OAI211_X1 g532(.A(new_n725_), .B(new_n529_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n727_), .A2(new_n330_), .A3(new_n529_), .A4(new_n724_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G99gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G99gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(G1338gat));
  XNOR2_X1  g540(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n727_), .A2(new_n330_), .A3(new_n634_), .A4(new_n724_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(G106gat), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n744_), .A2(new_n743_), .A3(G106gat), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n725_), .A2(new_n272_), .A3(new_n634_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n742_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n747_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n749_), .B(new_n742_), .C1(new_n751_), .C2(new_n745_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n750_), .A2(new_n753_), .ZN(G1339gat));
  NAND3_X1  g553(.A1(new_n664_), .A2(new_n610_), .A3(new_n693_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(KEYINPUT54), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(KEYINPUT54), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n755_), .A2(KEYINPUT54), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n311_), .A2(new_n316_), .A3(new_n313_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT55), .B(new_n316_), .C1(new_n311_), .C2(new_n313_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n325_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(new_n325_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n244_), .A4(new_n328_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n761_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n318_), .A2(KEYINPUT55), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n314_), .A2(new_n762_), .A3(new_n317_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n327_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n765_), .A2(new_n766_), .A3(new_n325_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n776_), .A2(new_n244_), .A3(new_n328_), .A4(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT114), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n230_), .A2(new_n231_), .A3(new_n221_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n218_), .A2(new_n220_), .A3(new_n232_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n240_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n243_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT115), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n771_), .A2(new_n779_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n640_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n783_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n776_), .A2(new_n328_), .A3(new_n777_), .A4(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT58), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(KEYINPUT116), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(KEYINPUT116), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n769_), .A2(new_n328_), .A3(new_n794_), .A4(new_n790_), .ZN(new_n795_));
  AND4_X1   g594(.A1(new_n577_), .A2(new_n793_), .A3(new_n795_), .A4(new_n583_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n786_), .A2(KEYINPUT57), .A3(new_n640_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n789_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n759_), .A2(new_n760_), .B1(new_n799_), .B2(new_n604_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n622_), .A2(new_n376_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n533_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G113gat), .B1(new_n803_), .B2(new_n244_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n786_), .A2(KEYINPUT57), .A3(new_n640_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT57), .B1(new_n786_), .B2(new_n640_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n796_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT117), .B1(new_n807_), .B2(new_n611_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n758_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n755_), .A2(new_n756_), .A3(KEYINPUT54), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n760_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n799_), .A2(new_n812_), .A3(new_n604_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n808_), .A2(new_n811_), .A3(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n802_), .A2(KEYINPUT59), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT59), .B1(new_n800_), .B2(new_n802_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n244_), .A2(G113gat), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n804_), .B1(new_n818_), .B2(new_n819_), .ZN(G1340gat));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n331_), .A3(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT118), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n816_), .A2(new_n823_), .A3(new_n817_), .A4(new_n331_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(G120gat), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT60), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n610_), .B2(G120gat), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n803_), .B(new_n827_), .C1(new_n826_), .C2(G120gat), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(G1341gat));
  AOI21_X1  g628(.A(G127gat), .B1(new_n803_), .B2(new_n611_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n611_), .A2(G127gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n818_), .B2(new_n831_), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(new_n803_), .B2(new_n570_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n584_), .A2(G134gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n818_), .B2(new_n834_), .ZN(G1343gat));
  NAND2_X1  g634(.A1(new_n799_), .A2(new_n604_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n801_), .A2(new_n535_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n811_), .A2(new_n836_), .B1(KEYINPUT119), .B2(new_n837_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n837_), .A2(KEYINPUT119), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n244_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g642(.A1(new_n840_), .A2(new_n332_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT120), .B(G148gat), .Z(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1345gat));
  NOR2_X1   g645(.A1(new_n840_), .A2(new_n604_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT61), .B(G155gat), .Z(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1346gat));
  AND3_X1   g648(.A1(new_n841_), .A2(G162gat), .A3(new_n584_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G162gat), .B1(new_n841_), .B2(new_n570_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1347gat));
  NOR2_X1   g651(.A1(new_n528_), .A2(new_n377_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n529_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n814_), .A2(new_n244_), .A3(new_n518_), .A4(new_n855_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n856_), .A2(G169gat), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n396_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT62), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(G169gat), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(G1348gat));
  NAND4_X1  g662(.A1(new_n814_), .A2(new_n330_), .A3(new_n518_), .A4(new_n855_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n393_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(KEYINPUT121), .A3(new_n393_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n800_), .A2(new_n634_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n332_), .A2(new_n393_), .A3(new_n854_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n867_), .A2(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1349gat));
  AND3_X1   g670(.A1(new_n814_), .A2(new_n518_), .A3(new_n855_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n604_), .A2(new_n415_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(new_n611_), .A3(new_n855_), .ZN(new_n874_));
  INV_X1    g673(.A(G183gat), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n872_), .A2(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1350gat));
  NAND3_X1  g675(.A1(new_n872_), .A2(new_n570_), .A3(new_n416_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n814_), .A2(new_n518_), .A3(new_n584_), .A4(new_n855_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n878_), .A2(new_n879_), .A3(G190gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n878_), .B2(G190gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n877_), .B1(new_n880_), .B2(new_n881_), .ZN(G1351gat));
  NOR2_X1   g681(.A1(new_n800_), .A2(new_n534_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n883_), .A2(new_n853_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(G197gat), .A4(new_n244_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n244_), .A3(new_n853_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n237_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT123), .B1(new_n887_), .B2(new_n237_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n886_), .A2(new_n888_), .A3(new_n889_), .ZN(G1352gat));
  AND3_X1   g689(.A1(new_n883_), .A2(new_n331_), .A3(new_n853_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT124), .B(G204gat), .Z(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n891_), .B2(new_n894_), .ZN(G1353gat));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n611_), .B1(new_n896_), .B2(new_n594_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT125), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n884_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n594_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1354gat));
  NAND2_X1  g700(.A1(new_n811_), .A2(new_n836_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n902_), .A2(new_n570_), .A3(new_n535_), .A4(new_n853_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT127), .B(G218gat), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n904_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n905_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n884_), .A2(new_n584_), .A3(new_n906_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1355gat));
endmodule


