//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT88), .B(G204gat), .Z(new_n209_));
  INV_X1    g008(.A(G197gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G204gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT21), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(G197gat), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n212_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT89), .B1(new_n212_), .B2(G197gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OAI221_X1 g016(.A(new_n208_), .B1(new_n211_), .B2(new_n213_), .C1(new_n217_), .C2(KEYINPUT21), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT21), .A3(new_n207_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT84), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n224_), .B2(new_n221_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n227_), .A2(KEYINPUT85), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(KEYINPUT85), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G169gat), .ZN(new_n232_));
  INV_X1    g031(.A(G176gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT26), .B(G190gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT25), .B(G183gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n228_), .A2(new_n229_), .A3(new_n234_), .A4(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(new_n224_), .B2(KEYINPUT23), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(G183gat), .B2(G190gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G169gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n220_), .B1(new_n238_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT20), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n218_), .A2(new_n219_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n236_), .B(KEYINPUT92), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n235_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n226_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n249_), .A2(new_n240_), .A3(new_n250_), .A4(new_n234_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n243_), .B1(new_n225_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n247_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT19), .ZN(new_n257_));
  NOR4_X1   g056(.A1(new_n245_), .A2(new_n246_), .A3(new_n255_), .A4(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n238_), .A2(new_n220_), .A3(new_n244_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n246_), .B1(new_n247_), .B2(new_n254_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n206_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n255_), .A2(new_n246_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n238_), .A2(new_n244_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n265_), .B1(new_n266_), .B2(new_n220_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n264_), .B(new_n205_), .C1(new_n267_), .C2(new_n257_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT27), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n271_), .A2(KEYINPUT101), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(KEYINPUT101), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n267_), .A2(new_n257_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT99), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n267_), .A2(KEYINPUT99), .A3(new_n257_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n260_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT100), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n280_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n277_), .A2(new_n278_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(new_n205_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n268_), .A2(KEYINPUT27), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n274_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT3), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT2), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT87), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n292_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(KEYINPUT1), .B2(new_n293_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(KEYINPUT1), .B2(new_n293_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n287_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(new_n289_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G127gat), .B(G134gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G113gat), .B(G120gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  NAND3_X1  g104(.A1(new_n301_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT95), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT96), .Z(new_n309_));
  AND2_X1   g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT94), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n301_), .A2(new_n305_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT93), .ZN(new_n313_));
  INV_X1    g112(.A(new_n305_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n296_), .A2(new_n300_), .A3(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n301_), .A2(KEYINPUT93), .A3(new_n305_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n311_), .B1(new_n318_), .B2(KEYINPUT4), .ZN(new_n319_));
  AOI211_X1 g118(.A(KEYINPUT94), .B(new_n302_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n310_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n308_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G1gat), .B(G29gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT97), .B(G85gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT0), .B(G57gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  NAND2_X1  g128(.A1(new_n324_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n329_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n321_), .A2(new_n323_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n220_), .B1(new_n301_), .B2(KEYINPUT29), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n335_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G78gat), .B(G106gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT90), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n338_), .B(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n301_), .A2(KEYINPUT29), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT28), .ZN(new_n343_));
  XOR2_X1   g142(.A(G22gat), .B(G50gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n336_), .A2(new_n337_), .A3(new_n340_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n347_), .A2(KEYINPUT91), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(KEYINPUT91), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n338_), .A2(new_n339_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n345_), .A2(new_n348_), .A3(new_n349_), .A4(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G15gat), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n266_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n266_), .A2(new_n354_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT31), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359_));
  INV_X1    g158(.A(G43gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(new_n305_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n358_), .B(new_n364_), .ZN(new_n365_));
  NOR4_X1   g164(.A1(new_n286_), .A2(new_n333_), .A3(new_n352_), .A4(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n264_), .B(new_n367_), .C1(new_n267_), .C2(new_n257_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n283_), .B2(new_n367_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n322_), .B(new_n306_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n331_), .B1(new_n318_), .B2(new_n309_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n269_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n321_), .A2(KEYINPUT33), .A3(new_n323_), .A4(new_n331_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT98), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n332_), .B2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n332_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n370_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n330_), .A2(new_n332_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n352_), .ZN(new_n383_));
  OAI22_X1  g182(.A1(new_n381_), .A2(new_n352_), .B1(new_n383_), .B2(new_n286_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n366_), .B1(new_n384_), .B2(new_n365_), .ZN(new_n385_));
  AND2_X1   g184(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G106gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G99gat), .A2(G106gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT6), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(G99gat), .A3(G106gat), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n388_), .A2(new_n389_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G85gat), .ZN(new_n395_));
  INV_X1    g194(.A(G92gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT9), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G85gat), .A2(G92gat), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n397_), .A2(KEYINPUT64), .A3(new_n398_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n397_), .ZN(new_n401_));
  AND2_X1   g200(.A1(G85gat), .A2(G92gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G85gat), .A2(G92gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n398_), .B1(new_n404_), .B2(KEYINPUT64), .ZN(new_n405_));
  OAI211_X1 g204(.A(KEYINPUT65), .B(new_n394_), .C1(new_n401_), .C2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n397_), .A2(KEYINPUT64), .A3(new_n399_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT9), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT65), .B1(new_n410_), .B2(new_n394_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n391_), .A2(new_n393_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT7), .ZN(new_n414_));
  INV_X1    g213(.A(G99gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n389_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n404_), .B1(new_n413_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT8), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n392_), .B1(G99gat), .B2(G106gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n390_), .A2(KEYINPUT6), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n417_), .B(new_n416_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT8), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n404_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G57gat), .B(G64gat), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT11), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(KEYINPUT11), .ZN(new_n429_));
  XOR2_X1   g228(.A(G71gat), .B(G78gat), .Z(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n429_), .A2(new_n430_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n412_), .A2(new_n426_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n412_), .A2(new_n426_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n433_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n437_), .B2(KEYINPUT66), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(KEYINPUT66), .B2(new_n437_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(G230gat), .A3(G233gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n397_), .A2(new_n399_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n417_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n391_), .A2(new_n393_), .ZN(new_n445_));
  AOI211_X1 g244(.A(KEYINPUT8), .B(new_n441_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n424_), .B1(new_n423_), .B2(new_n404_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT67), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n420_), .A2(new_n449_), .A3(new_n425_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n451_), .A2(KEYINPUT68), .A3(new_n412_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT68), .B1(new_n451_), .B2(new_n412_), .ZN(new_n453_));
  OAI211_X1 g252(.A(KEYINPUT12), .B(new_n436_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n434_), .B1(new_n437_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G230gat), .A2(G233gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n440_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G120gat), .B(G148gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT5), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G176gat), .B(G204gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n461_), .B(new_n462_), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n463_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n440_), .A2(new_n458_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT13), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n464_), .A2(KEYINPUT13), .A3(new_n466_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT15), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476_));
  INV_X1    g275(.A(G1gat), .ZN(new_n477_));
  INV_X1    g276(.A(G8gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n475_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n475_), .A2(KEYINPUT81), .A3(new_n482_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT80), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n474_), .A2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n474_), .A2(new_n487_), .ZN(new_n489_));
  OR3_X1    g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n482_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(new_n486_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT82), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OR3_X1    g293(.A1(new_n491_), .A2(KEYINPUT83), .A3(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT83), .B1(new_n491_), .B2(new_n494_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n482_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n490_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G229gat), .A3(G233gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(new_n496_), .A3(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G169gat), .B(G197gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n495_), .A2(new_n496_), .A3(new_n499_), .A4(new_n503_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n471_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n385_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G231gat), .A2(G233gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n433_), .B(new_n511_), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT77), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(new_n482_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G127gat), .B(G155gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(G183gat), .B(G211gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT17), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n519_), .A2(KEYINPUT17), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n514_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT79), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n522_), .B(KEYINPUT79), .C1(new_n514_), .C2(new_n520_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G190gat), .B(G218gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G134gat), .B(G162gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n529_), .B(KEYINPUT36), .Z(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n451_), .A2(new_n412_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n451_), .A2(new_n412_), .A3(KEYINPUT68), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT70), .B1(new_n536_), .B2(new_n475_), .ZN(new_n537_));
  OAI211_X1 g336(.A(KEYINPUT70), .B(new_n475_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT71), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n475_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT70), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT71), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n538_), .ZN(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n546_));
  NAND2_X1  g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(KEYINPUT35), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT72), .Z(new_n550_));
  NAND3_X1  g349(.A1(new_n412_), .A2(new_n474_), .A3(new_n426_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n540_), .A2(new_n545_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n548_), .A2(KEYINPUT35), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n555_), .B(KEYINPUT73), .ZN(new_n558_));
  AOI211_X1 g357(.A(new_n552_), .B(new_n558_), .C1(new_n543_), .C2(new_n538_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n531_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n529_), .A2(KEYINPUT36), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI211_X1 g362(.A(new_n563_), .B(new_n559_), .C1(new_n554_), .C2(new_n556_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT37), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT74), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n543_), .A2(new_n538_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n552_), .B1(new_n567_), .B2(KEYINPUT71), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n555_), .B1(new_n568_), .B2(new_n545_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n530_), .B1(new_n569_), .B2(new_n559_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n557_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT74), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(KEYINPUT37), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n566_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n559_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT75), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT75), .B1(new_n569_), .B2(new_n559_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n530_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n571_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n526_), .B1(new_n575_), .B2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n510_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n333_), .B(KEYINPUT102), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n477_), .A3(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT38), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n530_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n569_), .A2(KEYINPUT75), .A3(new_n559_), .ZN(new_n589_));
  OAI211_X1 g388(.A(KEYINPUT103), .B(new_n571_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT103), .B1(new_n580_), .B2(new_n571_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n525_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n510_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n596_), .B2(new_n382_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n587_), .A2(new_n597_), .ZN(G1324gat));
  NOR2_X1   g397(.A1(new_n284_), .A2(new_n285_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT104), .B1(new_n596_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n378_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n602_), .A2(new_n380_), .A3(new_n374_), .A4(new_n373_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n370_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n352_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n286_), .A2(new_n383_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n365_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n366_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n508_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n594_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n286_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT105), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n478_), .B1(new_n614_), .B2(KEYINPUT39), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n601_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n614_), .A2(KEYINPUT39), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n601_), .A2(new_n613_), .A3(new_n615_), .A4(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n584_), .A2(new_n478_), .A3(new_n286_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n618_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n618_), .A2(new_n620_), .A3(KEYINPUT40), .A4(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1325gat));
  INV_X1    g425(.A(G15gat), .ZN(new_n627_));
  INV_X1    g426(.A(new_n365_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n611_), .B2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT41), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n584_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1326gat));
  INV_X1    g431(.A(new_n352_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G22gat), .B1(new_n596_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n584_), .A2(new_n636_), .A3(new_n352_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1327gat));
  NOR2_X1   g437(.A1(new_n593_), .A2(new_n525_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n510_), .A2(new_n639_), .ZN(new_n640_));
  OR3_X1    g439(.A1(new_n640_), .A2(G29gat), .A3(new_n382_), .ZN(new_n641_));
  OR2_X1    g440(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n642_));
  NAND2_X1  g441(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n573_), .B1(new_n572_), .B2(KEYINPUT37), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT37), .ZN(new_n645_));
  AOI211_X1 g444(.A(KEYINPUT74), .B(new_n645_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n582_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n642_), .B(new_n643_), .C1(new_n385_), .C2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n647_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n609_), .A2(KEYINPUT106), .A3(KEYINPUT43), .A4(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n509_), .A2(new_n525_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n648_), .A2(new_n650_), .A3(KEYINPUT44), .A4(new_n651_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n585_), .A3(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n656_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT107), .B1(new_n656_), .B2(G29gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n641_), .B1(new_n657_), .B2(new_n658_), .ZN(G1328gat));
  NOR3_X1   g458(.A1(new_n640_), .A2(G36gat), .A3(new_n600_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT45), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n654_), .A2(new_n286_), .A3(new_n655_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G36gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(new_n664_), .A3(KEYINPUT46), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  NAND4_X1  g468(.A1(new_n654_), .A2(G43gat), .A3(new_n628_), .A4(new_n655_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n360_), .B1(new_n640_), .B2(new_n365_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g472(.A1(new_n640_), .A2(G50gat), .A3(new_n633_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n654_), .A2(new_n352_), .A3(new_n655_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(new_n676_), .A3(G50gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n675_), .B2(G50gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(G1331gat));
  INV_X1    g478(.A(new_n471_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n507_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n385_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n595_), .ZN(new_n685_));
  INV_X1    g484(.A(G57gat), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(new_n382_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n585_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n684_), .A2(new_n583_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n691_), .B1(new_n690_), .B2(new_n689_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n686_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n692_), .A2(KEYINPUT110), .A3(new_n686_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n687_), .B1(new_n695_), .B2(new_n696_), .ZN(G1332gat));
  OAI21_X1  g496(.A(G64gat), .B1(new_n685_), .B2(new_n600_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT48), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n600_), .A2(G64gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n689_), .B2(new_n700_), .ZN(G1333gat));
  OAI21_X1  g500(.A(G71gat), .B1(new_n685_), .B2(new_n365_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT49), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n365_), .A2(G71gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n689_), .B2(new_n704_), .ZN(G1334gat));
  OAI21_X1  g504(.A(G78gat), .B1(new_n685_), .B2(new_n633_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT50), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n633_), .A2(G78gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n689_), .B2(new_n708_), .ZN(G1335gat));
  NOR2_X1   g508(.A1(new_n683_), .A2(new_n525_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n648_), .A2(new_n650_), .A3(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n382_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n684_), .A2(new_n639_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n395_), .A3(new_n585_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1336gat));
  OAI21_X1  g514(.A(G92gat), .B1(new_n711_), .B2(new_n600_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n713_), .A2(new_n396_), .A3(new_n286_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT111), .ZN(G1337gat));
  OAI21_X1  g518(.A(G99gat), .B1(new_n711_), .B2(new_n365_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n713_), .A2(new_n388_), .A3(new_n628_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g522(.A1(new_n713_), .A2(new_n389_), .A3(new_n352_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n648_), .A2(new_n650_), .A3(new_n352_), .A4(new_n710_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(G106gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(G106gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g529(.A(KEYINPUT115), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n471_), .A2(new_n681_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n583_), .B2(new_n734_), .ZN(new_n735_));
  AND4_X1   g534(.A1(new_n525_), .A2(new_n647_), .A3(new_n733_), .A4(new_n734_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n571_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n457_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n458_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n454_), .A2(new_n456_), .A3(KEYINPUT55), .A4(new_n457_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT56), .B1(new_n745_), .B2(new_n463_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  AOI211_X1 g546(.A(new_n747_), .B(new_n465_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n681_), .B(new_n466_), .C1(new_n746_), .C2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n503_), .B1(new_n498_), .B2(new_n493_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(new_n493_), .B2(new_n491_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n506_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n467_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n749_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(KEYINPUT57), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n740_), .A2(new_n590_), .A3(new_n754_), .A4(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n746_), .A2(new_n748_), .A3(KEYINPUT114), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n745_), .A2(new_n463_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(KEYINPUT114), .A3(new_n747_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n752_), .A2(new_n466_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n759_), .B1(new_n760_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n746_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n745_), .A2(KEYINPUT56), .A3(new_n463_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n769_), .A2(KEYINPUT58), .A3(new_n762_), .A4(new_n763_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n765_), .A2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n758_), .B1(new_n647_), .B2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n757_), .B1(new_n593_), .B2(new_n754_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n526_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n737_), .A2(new_n774_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n286_), .A2(new_n352_), .A3(new_n365_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n585_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n731_), .B1(new_n775_), .B2(new_n778_), .ZN(new_n779_));
  AOI211_X1 g578(.A(KEYINPUT115), .B(new_n777_), .C1(new_n737_), .C2(new_n774_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G113gat), .B1(new_n781_), .B2(new_n681_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT59), .B1(new_n775_), .B2(new_n778_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT59), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n785_), .B(new_n777_), .C1(new_n737_), .C2(new_n774_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n647_), .A2(new_n771_), .ZN(new_n788_));
  AND4_X1   g587(.A1(new_n740_), .A2(new_n590_), .A3(new_n754_), .A4(new_n757_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n593_), .A2(new_n754_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n756_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n525_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n583_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n647_), .A2(new_n525_), .A3(new_n734_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n732_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n778_), .B1(new_n793_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n785_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n777_), .B1(new_n737_), .B2(new_n774_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT59), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(KEYINPUT116), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n787_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(G113gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n681_), .B2(KEYINPUT117), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(KEYINPUT117), .B2(new_n804_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n782_), .B1(new_n803_), .B2(new_n806_), .ZN(G1340gat));
  AOI21_X1  g606(.A(new_n680_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n808_));
  INV_X1    g607(.A(G120gat), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n798_), .A2(KEYINPUT115), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n800_), .A2(new_n731_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n809_), .B1(new_n680_), .B2(KEYINPUT60), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(KEYINPUT60), .B2(new_n809_), .ZN(new_n814_));
  OAI22_X1  g613(.A1(new_n808_), .A2(new_n809_), .B1(new_n812_), .B2(new_n814_), .ZN(G1341gat));
  INV_X1    g614(.A(G127gat), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n526_), .A2(new_n816_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n784_), .A2(new_n786_), .A3(new_n783_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT116), .B1(new_n799_), .B2(new_n801_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n812_), .B2(new_n526_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(KEYINPUT118), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823_));
  INV_X1    g622(.A(new_n817_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n787_), .B2(new_n802_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G127gat), .B1(new_n781_), .B2(new_n525_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n823_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n822_), .A2(new_n827_), .ZN(G1342gat));
  NAND3_X1  g627(.A1(new_n803_), .A2(G134gat), .A3(new_n649_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n593_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n810_), .A2(new_n830_), .A3(new_n811_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832_));
  INV_X1    g631(.A(G134gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n833_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT119), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n829_), .A2(new_n834_), .A3(new_n836_), .ZN(G1343gat));
  NOR4_X1   g636(.A1(new_n688_), .A2(new_n633_), .A3(new_n286_), .A4(new_n628_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n775_), .A2(new_n838_), .ZN(new_n839_));
  OR3_X1    g638(.A1(new_n839_), .A2(KEYINPUT121), .A3(new_n507_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT121), .B1(new_n839_), .B2(new_n507_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT120), .B(G141gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1344gat));
  INV_X1    g643(.A(new_n839_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n471_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g646(.A1(new_n839_), .A2(new_n526_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT61), .B(G155gat), .Z(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  OR3_X1    g649(.A1(new_n839_), .A2(G162gat), .A3(new_n593_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G162gat), .B1(new_n839_), .B2(new_n647_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1347gat));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n585_), .A2(new_n600_), .A3(new_n365_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n775_), .A2(new_n633_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n681_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n854_), .B1(new_n858_), .B2(G169gat), .ZN(new_n859_));
  AOI211_X1 g658(.A(KEYINPUT62), .B(new_n232_), .C1(new_n857_), .C2(new_n681_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n856_), .A2(KEYINPUT122), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n775_), .A2(new_n862_), .A3(new_n633_), .A4(new_n855_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n866_));
  AND2_X1   g665(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n681_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n859_), .A2(new_n860_), .B1(new_n865_), .B2(new_n868_), .ZN(G1348gat));
  INV_X1    g668(.A(new_n855_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n775_), .A2(new_n633_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT123), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n775_), .A2(new_n873_), .A3(new_n633_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n870_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n680_), .A2(new_n233_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n875_), .B2(new_n877_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G176gat), .B1(new_n864_), .B2(new_n471_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(G1349gat));
  NOR2_X1   g680(.A1(new_n526_), .A2(new_n248_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n864_), .A2(KEYINPUT125), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(G183gat), .B1(new_n875_), .B2(new_n525_), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT125), .B1(new_n864_), .B2(new_n882_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n865_), .B2(new_n647_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n864_), .A2(new_n235_), .A3(new_n830_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1351gat));
  NOR3_X1   g688(.A1(new_n383_), .A2(new_n600_), .A3(new_n628_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n775_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n681_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n471_), .ZN(new_n894_));
  MUX2_X1   g693(.A(new_n209_), .B(G204gat), .S(new_n894_), .Z(G1353gat));
  AOI21_X1  g694(.A(new_n526_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n891_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT126), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n891_), .A2(new_n899_), .A3(new_n896_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1354gat));
  INV_X1    g702(.A(new_n891_), .ZN(new_n904_));
  OR3_X1    g703(.A1(new_n904_), .A2(G218gat), .A3(new_n593_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G218gat), .B1(new_n904_), .B2(new_n647_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1355gat));
endmodule


