//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n978_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n985_, new_n986_, new_n987_;
  NOR2_X1   g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n205_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT66), .B1(new_n207_), .B2(new_n202_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI22_X1  g012(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n213_), .B(new_n214_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n209_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(new_n209_), .B2(new_n218_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n203_), .A2(KEYINPUT9), .A3(new_n205_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT10), .B(G99gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT64), .B(G85gat), .ZN(new_n225_));
  INV_X1    g024(.A(G92gat), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(KEYINPUT9), .ZN(new_n227_));
  OAI22_X1  g026(.A1(G106gat), .A2(new_n224_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  OAI22_X1  g027(.A1(new_n220_), .A2(new_n221_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G57gat), .B(G64gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G78gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT11), .ZN(new_n232_));
  XOR2_X1   g031(.A(G71gat), .B(G78gat), .Z(new_n233_));
  INV_X1    g032(.A(G64gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G57gat), .ZN(new_n235_));
  INV_X1    g034(.A(G57gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G64gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n237_), .A3(KEYINPUT11), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n232_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT67), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n243_), .B(new_n232_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n229_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT12), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G230gat), .A2(G233gat), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n242_), .A2(new_n244_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n223_), .A2(new_n228_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n209_), .A2(new_n218_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT8), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n209_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n251_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n241_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n229_), .A2(KEYINPUT12), .A3(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n248_), .A2(new_n249_), .A3(new_n256_), .A4(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n246_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n249_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT12), .B(new_n232_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n255_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n229_), .A2(new_n245_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n268_), .A2(KEYINPUT68), .A3(new_n249_), .A4(new_n248_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n261_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT5), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G176gat), .B(G204gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n261_), .A2(new_n264_), .A3(new_n269_), .A4(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT13), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT69), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT13), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n278_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G29gat), .B(G36gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G43gat), .B(G50gat), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT70), .B(KEYINPUT15), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n229_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n255_), .A2(new_n290_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G232gat), .A2(G233gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT34), .Z(new_n296_));
  INV_X1    g095(.A(KEYINPUT35), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT71), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n296_), .A2(new_n297_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n293_), .A2(new_n294_), .A3(new_n299_), .A4(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n300_), .A2(new_n301_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n303_), .A2(new_n304_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G190gat), .B(G218gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT72), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G134gat), .B(G162gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT36), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n311_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n314_), .A2(KEYINPUT36), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT37), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT37), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n313_), .A2(new_n319_), .A3(new_n316_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G15gat), .B(G22gat), .ZN(new_n323_));
  INV_X1    g122(.A(G1gat), .ZN(new_n324_));
  INV_X1    g123(.A(G8gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT14), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G1gat), .B(G8gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G231gat), .A2(G233gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT76), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n332_), .A2(new_n250_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n250_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G127gat), .B(G155gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G183gat), .B(G211gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT17), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT77), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n333_), .A2(new_n334_), .A3(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n331_), .B(KEYINPUT74), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n343_), .A2(new_n257_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n257_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT17), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n339_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n342_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n322_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n285_), .A2(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n351_), .B(KEYINPUT78), .Z(new_n352_));
  NAND2_X1  g151(.A1(G228gat), .A2(G233gat), .ZN(new_n353_));
  INV_X1    g152(.A(G218gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G211gat), .ZN(new_n355_));
  INV_X1    g154(.A(G211gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G218gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G204gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G197gat), .ZN(new_n360_));
  INV_X1    g159(.A(G197gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(G204gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n358_), .B1(KEYINPUT21), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(KEYINPUT89), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n359_), .A3(G197gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT21), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n365_), .A2(new_n367_), .A3(new_n368_), .A4(new_n362_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n367_), .A3(new_n362_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n353_), .B1(new_n374_), .B2(KEYINPUT90), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G155gat), .A2(G162gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT86), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(G155gat), .A3(G162gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT87), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n384_), .B(new_n390_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  AOI211_X1 g192(.A(KEYINPUT87), .B(new_n389_), .C1(new_n386_), .C2(new_n388_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n383_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT88), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n382_), .B(KEYINPUT3), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n397_), .B(new_n398_), .C1(KEYINPUT2), .C2(new_n381_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n386_), .A2(new_n388_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n384_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n376_), .B1(new_n395_), .B2(new_n403_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n364_), .A2(new_n369_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n405_));
  OAI21_X1  g204(.A(G78gat), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G78gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(KEYINPUT1), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT87), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n390_), .A2(new_n384_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n391_), .A2(new_n392_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n412_), .A2(new_n383_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n407_), .B(new_n374_), .C1(new_n413_), .C2(new_n376_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n406_), .A2(new_n414_), .A3(G106gat), .ZN(new_n415_));
  AOI21_X1  g214(.A(G106gat), .B1(new_n406_), .B2(new_n414_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n375_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n381_), .A2(new_n382_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n392_), .B1(new_n400_), .B2(KEYINPUT1), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n390_), .A2(new_n384_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(new_n421_), .B2(new_n411_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT3), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n382_), .B(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT2), .B1(new_n379_), .B2(new_n380_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n401_), .B1(new_n426_), .B2(new_n397_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT29), .B1(new_n422_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n407_), .B1(new_n428_), .B2(new_n374_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n404_), .A2(G78gat), .A3(new_n405_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n212_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n406_), .A2(new_n414_), .A3(G106gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n375_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n395_), .A2(new_n403_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT28), .B1(new_n435_), .B2(KEYINPUT29), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT28), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n413_), .A2(new_n437_), .A3(new_n376_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G22gat), .B(G50gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n436_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n417_), .A2(new_n434_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n417_), .B2(new_n434_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT93), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G127gat), .B(G134gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G113gat), .B(G120gat), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n450_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI211_X1 g252(.A(new_n448_), .B(new_n453_), .C1(new_n395_), .C2(new_n403_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n452_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT93), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n457_));
  AND4_X1   g256(.A1(new_n456_), .A2(new_n395_), .A3(new_n457_), .A4(new_n403_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n447_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G57gat), .B(G85gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT4), .ZN(new_n466_));
  OAI211_X1 g265(.A(KEYINPUT93), .B(new_n455_), .C1(new_n422_), .C2(new_n427_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n395_), .A2(new_n403_), .A3(new_n456_), .A4(new_n457_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT94), .B(KEYINPUT4), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n435_), .A2(new_n453_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n447_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n459_), .B(new_n465_), .C1(new_n469_), .C2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT4), .B1(new_n454_), .B2(new_n458_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n471_), .A2(new_n472_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n474_), .B1(new_n478_), .B2(new_n465_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT100), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n469_), .A2(new_n473_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n464_), .B1(new_n481_), .B2(new_n475_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT100), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n483_), .A3(new_n474_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n446_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT27), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G8gat), .B(G36gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G64gat), .B(G92gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(G169gat), .A2(G176gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(KEYINPUT24), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT25), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT79), .B1(new_n497_), .B2(G183gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT79), .ZN(new_n499_));
  INV_X1    g298(.A(G183gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT25), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(G183gat), .ZN(new_n503_));
  INV_X1    g302(.A(G190gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT26), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT26), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G190gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n503_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n496_), .B1(new_n502_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT80), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT80), .B(new_n496_), .C1(new_n502_), .C2(new_n508_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n494_), .A2(KEYINPUT24), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G183gat), .A2(G190gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT23), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT81), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n514_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT23), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(G183gat), .A3(G190gat), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n513_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n511_), .A2(new_n512_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n515_), .A2(new_n521_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(G183gat), .B2(G190gat), .ZN(new_n525_));
  INV_X1    g324(.A(G176gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT22), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n526_), .B1(new_n527_), .B2(KEYINPUT82), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(G169gat), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n528_), .A2(G169gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n525_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n405_), .B1(new_n523_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n495_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G169gat), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n534_), .B2(new_n526_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n521_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n536_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(G183gat), .A2(G190gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n535_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT26), .B(G190gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n500_), .A2(KEYINPUT25), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(new_n503_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n513_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n496_), .A4(new_n524_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n405_), .A2(new_n539_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G226gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT19), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n532_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n539_), .A2(new_n544_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n552_), .B2(new_n374_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n522_), .A2(new_n512_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n540_), .A2(new_n503_), .A3(new_n498_), .A4(new_n501_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT80), .B1(new_n555_), .B2(new_n496_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n405_), .B(new_n531_), .C1(new_n554_), .C2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n551_), .A2(KEYINPUT91), .B1(new_n558_), .B2(new_n547_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n532_), .B2(new_n550_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n493_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n547_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n531_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n374_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n565_), .A2(KEYINPUT91), .A3(new_n545_), .A4(new_n549_), .ZN(new_n566_));
  AND4_X1   g365(.A1(new_n493_), .A2(new_n563_), .A3(new_n566_), .A4(new_n561_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n487_), .B1(new_n562_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT102), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT102), .B(new_n487_), .C1(new_n562_), .C2(new_n567_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n547_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n553_), .A2(new_n572_), .A3(new_n557_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n553_), .A2(new_n557_), .A3(KEYINPUT98), .A4(new_n572_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n545_), .A2(KEYINPUT20), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n547_), .B1(new_n532_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n579_), .A2(new_n492_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n563_), .A2(new_n566_), .A3(new_n493_), .A4(new_n561_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT27), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT101), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n492_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT101), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(KEYINPUT27), .A4(new_n581_), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n570_), .A2(new_n571_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n493_), .A2(KEYINPUT32), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n579_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT99), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n563_), .A2(new_n566_), .A3(new_n561_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(new_n588_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n579_), .A2(new_n593_), .A3(new_n588_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n590_), .A2(new_n479_), .A3(new_n592_), .A4(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n476_), .A2(new_n477_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n467_), .A2(new_n468_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n464_), .B1(new_n597_), .B2(new_n447_), .ZN(new_n598_));
  AOI211_X1 g397(.A(KEYINPUT96), .B(KEYINPUT33), .C1(new_n596_), .C2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n474_), .B2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n597_), .A2(new_n472_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT97), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n464_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n476_), .A2(new_n447_), .A3(new_n471_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n447_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT97), .B1(new_n608_), .B2(new_n465_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n606_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n591_), .A2(new_n492_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n596_), .A2(KEYINPUT33), .A3(new_n598_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n610_), .A2(new_n581_), .A3(new_n611_), .A4(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n595_), .B1(new_n603_), .B2(new_n613_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n486_), .A2(new_n587_), .B1(new_n614_), .B2(new_n446_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G71gat), .B(G99gat), .ZN(new_n616_));
  INV_X1    g415(.A(G43gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n564_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G227gat), .A2(G233gat), .ZN(new_n620_));
  INV_X1    g419(.A(G15gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT30), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT83), .ZN(new_n624_));
  INV_X1    g423(.A(new_n618_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n523_), .A2(new_n531_), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n619_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n624_), .B1(new_n619_), .B2(new_n626_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n628_), .A2(new_n629_), .A3(KEYINPUT31), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT31), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n619_), .A2(new_n626_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT83), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n623_), .B(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n631_), .B1(new_n635_), .B2(new_n627_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n455_), .B1(new_n630_), .B2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT31), .B1(new_n628_), .B2(new_n629_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n635_), .A2(new_n631_), .A3(new_n627_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n453_), .A3(new_n639_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n637_), .A2(KEYINPUT84), .A3(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT84), .B1(new_n637_), .B2(new_n640_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT103), .B1(new_n615_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n570_), .A2(new_n571_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n479_), .A2(KEYINPUT100), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n483_), .B1(new_n482_), .B2(new_n474_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n417_), .A2(new_n434_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n443_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n417_), .A2(new_n434_), .A3(new_n443_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n583_), .A2(new_n586_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n645_), .A2(new_n648_), .A3(new_n653_), .A4(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n614_), .A2(new_n446_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n658_));
  INV_X1    g457(.A(new_n643_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n637_), .A2(new_n640_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n587_), .A2(new_n648_), .A3(new_n446_), .A4(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n644_), .A2(new_n660_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n292_), .A2(new_n329_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n290_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n665_), .A2(new_n329_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(G229gat), .A2(G233gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n665_), .B(new_n329_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n667_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n668_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(G113gat), .B(G141gat), .ZN(new_n673_));
  XNOR2_X1  g472(.A(G169gat), .B(G197gat), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n673_), .B(new_n674_), .Z(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n672_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n668_), .A2(new_n671_), .A3(new_n675_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n663_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n352_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n324_), .A3(new_n485_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n663_), .A2(new_n317_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n280_), .A2(new_n284_), .A3(new_n679_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT104), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n280_), .A2(new_n284_), .A3(new_n686_), .A4(new_n679_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n683_), .A2(new_n688_), .A3(new_n349_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(new_n485_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n682_), .B1(new_n690_), .B2(new_n324_), .ZN(new_n691_));
  MUX2_X1   g490(.A(new_n682_), .B(new_n691_), .S(KEYINPUT38), .Z(G1324gat));
  INV_X1    g491(.A(new_n587_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n681_), .A2(new_n325_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(new_n693_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n325_), .B1(KEYINPUT105), .B2(KEYINPUT39), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT40), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(G1325gat));
  AOI21_X1  g501(.A(new_n621_), .B1(new_n689_), .B2(new_n643_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT41), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n681_), .A2(new_n621_), .A3(new_n643_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1326gat));
  INV_X1    g505(.A(G22gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n681_), .A2(new_n707_), .A3(new_n653_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n689_), .B2(new_n653_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n709_), .A2(new_n710_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(G1327gat));
  INV_X1    g512(.A(new_n285_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n317_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n349_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT107), .Z(new_n717_));
  NOR2_X1   g516(.A1(new_n714_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n680_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G29gat), .B1(new_n720_), .B2(new_n485_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n685_), .A2(new_n687_), .A3(new_n349_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n643_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n662_), .B1(new_n724_), .B2(new_n658_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n615_), .A2(KEYINPUT103), .A3(new_n643_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n723_), .B(new_n322_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n723_), .B1(new_n663_), .B2(new_n322_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n722_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n322_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT43), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n727_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(KEYINPUT44), .A3(new_n722_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n732_), .A2(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n485_), .A2(G29gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n721_), .B1(new_n737_), .B2(new_n738_), .ZN(G1328gat));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n587_), .A2(G36gat), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n719_), .B2(new_n742_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n680_), .A2(KEYINPUT45), .A3(new_n718_), .A4(new_n741_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n732_), .A2(new_n693_), .A3(new_n736_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(G36gat), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n748_), .A2(new_n749_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n747_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n750_), .A2(new_n753_), .ZN(G1329gat));
  OAI21_X1  g553(.A(new_n617_), .B1(new_n719_), .B2(new_n659_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT109), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n732_), .A2(new_n736_), .A3(G43gat), .A4(new_n661_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT47), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(new_n760_), .A3(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1330gat));
  AOI21_X1  g561(.A(G50gat), .B1(new_n720_), .B2(new_n653_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n653_), .A2(G50gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n737_), .B2(new_n764_), .ZN(G1331gat));
  INV_X1    g564(.A(new_n679_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n342_), .A2(new_n348_), .A3(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n285_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n663_), .A3(new_n317_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G57gat), .B1(new_n769_), .B2(new_n648_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n663_), .A2(new_n766_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n285_), .A2(new_n349_), .A3(new_n322_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n485_), .A2(new_n236_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1332gat));
  OAI21_X1  g574(.A(G64gat), .B1(new_n769_), .B2(new_n587_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT48), .ZN(new_n777_));
  INV_X1    g576(.A(new_n773_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n234_), .A3(new_n693_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT110), .ZN(G1333gat));
  OAI21_X1  g580(.A(G71gat), .B1(new_n769_), .B2(new_n659_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT49), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n659_), .A2(G71gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n773_), .B2(new_n784_), .ZN(G1334gat));
  NAND3_X1  g584(.A1(new_n778_), .A2(new_n407_), .A3(new_n653_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G78gat), .B1(new_n769_), .B2(new_n446_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT112), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n789_), .B(G78gat), .C1(new_n769_), .C2(new_n446_), .ZN(new_n790_));
  XOR2_X1   g589(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n791_));
  AND3_X1   g590(.A1(new_n788_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n786_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT113), .ZN(G1335gat));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n714_), .A2(new_n766_), .A3(new_n349_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n735_), .B2(new_n799_), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT114), .B(new_n798_), .C1(new_n734_), .C2(new_n727_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n796_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n799_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT114), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n735_), .A2(new_n797_), .A3(new_n799_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(KEYINPUT115), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n802_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n648_), .A2(new_n225_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(G85gat), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n285_), .A2(new_n717_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n771_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n812_), .B2(new_n648_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n809_), .A2(KEYINPUT116), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  INV_X1    g614(.A(new_n808_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n802_), .B2(new_n806_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n813_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n815_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n814_), .A2(new_n819_), .ZN(G1336gat));
  INV_X1    g619(.A(new_n812_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(new_n226_), .A3(new_n693_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n587_), .B1(new_n802_), .B2(new_n806_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n226_), .ZN(G1337gat));
  AOI21_X1  g623(.A(new_n659_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n661_), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n826_), .A2(new_n224_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n825_), .A2(new_n211_), .B1(new_n812_), .B2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g628(.A1(new_n821_), .A2(new_n212_), .A3(new_n653_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n735_), .A2(new_n653_), .A3(new_n799_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n831_), .A2(new_n832_), .A3(G106gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n831_), .B2(G106gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n830_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n693_), .A2(new_n653_), .A3(new_n826_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n349_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n675_), .B1(new_n669_), .B2(new_n667_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n664_), .A2(new_n666_), .A3(new_n670_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n678_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n278_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n256_), .A2(new_n258_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT12), .B1(new_n229_), .B2(new_n245_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847_));
  NOR4_X1   g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .A4(new_n263_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n249_), .B1(new_n268_), .B2(new_n248_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n261_), .A2(new_n847_), .A3(new_n269_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT56), .B1(new_n852_), .B2(new_n274_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n854_), .B(new_n276_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n277_), .A2(new_n679_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n277_), .A2(KEYINPUT117), .A3(new_n679_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n844_), .B1(new_n856_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n317_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n852_), .A2(new_n274_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n854_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n852_), .A2(KEYINPUT56), .A3(new_n274_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n277_), .B2(new_n843_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n277_), .A2(new_n869_), .A3(new_n843_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n868_), .B(KEYINPUT58), .C1(new_n870_), .C2(new_n871_), .ZN(new_n872_));
  OAI22_X1  g671(.A1(new_n853_), .A2(new_n855_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n321_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n863_), .A2(new_n864_), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n862_), .A2(KEYINPUT57), .A3(new_n317_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n839_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n767_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n279_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n279_), .B2(new_n879_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n485_), .B(new_n838_), .C1(new_n878_), .C2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT120), .B1(new_n878_), .B2(new_n883_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n844_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n861_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n868_), .B2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n864_), .B1(new_n890_), .B2(new_n715_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n875_), .A2(new_n872_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n877_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n883_), .B1(new_n893_), .B2(new_n349_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n838_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n894_), .A2(new_n648_), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n885_), .B1(new_n894_), .B2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n887_), .A2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n837_), .B1(new_n900_), .B2(new_n679_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n896_), .A2(KEYINPUT119), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n884_), .A2(new_n903_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n902_), .A2(new_n904_), .A3(new_n837_), .A4(new_n679_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT121), .B1(new_n901_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n766_), .B1(new_n887_), .B2(new_n899_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n908_), .B(new_n905_), .C1(new_n909_), .C2(new_n837_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n907_), .A2(new_n910_), .ZN(G1340gat));
  INV_X1    g710(.A(new_n900_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G120gat), .B1(new_n912_), .B2(new_n285_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n902_), .A2(new_n904_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n916_));
  AOI21_X1  g715(.A(G120gat), .B1(new_n714_), .B2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n916_), .B2(G120gat), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n914_), .A2(new_n915_), .A3(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n915_), .B1(new_n914_), .B2(new_n918_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n913_), .B1(new_n919_), .B2(new_n920_), .ZN(G1341gat));
  AOI21_X1  g720(.A(G127gat), .B1(new_n914_), .B2(new_n839_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n839_), .A2(G127gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT123), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n900_), .B2(new_n924_), .ZN(G1342gat));
  XOR2_X1   g724(.A(KEYINPUT124), .B(G134gat), .Z(new_n926_));
  NOR3_X1   g725(.A1(new_n912_), .A2(new_n321_), .A3(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(G134gat), .B1(new_n914_), .B2(new_n715_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1343gat));
  OAI21_X1  g728(.A(new_n485_), .B1(new_n878_), .B2(new_n883_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n659_), .A2(new_n653_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n930_), .A2(new_n693_), .A3(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n679_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n714_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g735(.A1(new_n932_), .A2(new_n839_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT61), .B(G155gat), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n937_), .B(new_n938_), .ZN(G1346gat));
  INV_X1    g738(.A(new_n932_), .ZN(new_n940_));
  OR3_X1    g739(.A1(new_n940_), .A2(G162gat), .A3(new_n317_), .ZN(new_n941_));
  OAI21_X1  g740(.A(G162gat), .B1(new_n940_), .B2(new_n321_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1347gat));
  NOR2_X1   g742(.A1(new_n587_), .A2(new_n485_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n894_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n659_), .A2(new_n653_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n946_), .A2(KEYINPUT125), .A3(new_n947_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n952_), .A2(new_n534_), .A3(new_n679_), .ZN(new_n953_));
  OAI21_X1  g752(.A(G169gat), .B1(new_n948_), .B2(new_n766_), .ZN(new_n954_));
  AND2_X1   g753(.A1(new_n954_), .A2(KEYINPUT62), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n954_), .A2(KEYINPUT62), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n953_), .B1(new_n955_), .B2(new_n956_), .ZN(G1348gat));
  NAND3_X1  g756(.A1(new_n952_), .A2(new_n526_), .A3(new_n714_), .ZN(new_n958_));
  OAI21_X1  g757(.A(G176gat), .B1(new_n948_), .B2(new_n285_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1349gat));
  NOR3_X1   g759(.A1(new_n948_), .A2(KEYINPUT126), .A3(new_n349_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(G183gat), .ZN(new_n962_));
  OAI21_X1  g761(.A(KEYINPUT126), .B1(new_n948_), .B2(new_n349_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n349_), .B1(new_n503_), .B2(new_n541_), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n962_), .A2(new_n963_), .B1(new_n952_), .B2(new_n964_), .ZN(G1350gat));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n504_), .B1(new_n952_), .B2(new_n322_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n715_), .A2(new_n540_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n968_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n966_), .B1(new_n967_), .B2(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n969_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n321_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n972_));
  OAI211_X1 g771(.A(new_n971_), .B(KEYINPUT127), .C1(new_n504_), .C2(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n970_), .A2(new_n973_), .ZN(G1351gat));
  NOR3_X1   g773(.A1(new_n894_), .A2(new_n931_), .A3(new_n945_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(new_n679_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n714_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g778(.A1(new_n975_), .A2(new_n839_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n981_));
  AND2_X1   g780(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n980_), .A2(new_n981_), .A3(new_n982_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n983_), .B1(new_n980_), .B2(new_n981_), .ZN(G1354gat));
  INV_X1    g783(.A(new_n975_), .ZN(new_n985_));
  OAI21_X1  g784(.A(G218gat), .B1(new_n985_), .B2(new_n321_), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n975_), .A2(new_n354_), .A3(new_n715_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n986_), .A2(new_n987_), .ZN(G1355gat));
endmodule


