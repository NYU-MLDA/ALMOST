//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT83), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT84), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n210_), .B2(KEYINPUT1), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT84), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n209_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n202_), .B(new_n205_), .C1(new_n211_), .C2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n205_), .A2(KEYINPUT3), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n202_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n205_), .A2(KEYINPUT3), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n210_), .A3(new_n208_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n216_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G120gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n227_), .B1(new_n216_), .B2(new_n223_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G225gat), .A2(G233gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(new_n232_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n229_), .A2(new_n234_), .A3(new_n230_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n233_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G1gat), .B(G29gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT0), .ZN(new_n240_));
  INV_X1    g039(.A(G57gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G85gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(new_n244_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n233_), .B(new_n243_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G78gat), .B(G106gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT28), .B1(new_n224_), .B2(KEYINPUT29), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n224_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n252_));
  XOR2_X1   g051(.A(G22gat), .B(G50gat), .Z(new_n253_));
  NOR3_X1   g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n252_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(new_n250_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n249_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT21), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G211gat), .B(G218gat), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n262_), .A2(KEYINPUT87), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(KEYINPUT87), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT86), .B(new_n261_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n259_), .A2(new_n260_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n265_), .B(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n268_), .B1(KEYINPUT29), .B2(new_n224_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G228gat), .A2(G233gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n270_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n269_), .B(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n253_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n256_), .A2(new_n250_), .A3(new_n255_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n249_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n274_), .B(new_n275_), .C1(KEYINPUT88), .C2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n258_), .A2(new_n273_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n273_), .B1(new_n258_), .B2(new_n277_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281_));
  INV_X1    g080(.A(G43gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G15gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n283_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT23), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(G183gat), .B2(G190gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT22), .B(G169gat), .ZN(new_n292_));
  INV_X1    g091(.A(G176gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n289_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT25), .B(G183gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT26), .B(G190gat), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n290_), .A2(KEYINPUT24), .ZN(new_n298_));
  OR2_X1    g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n296_), .A2(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n299_), .A2(KEYINPUT24), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n288_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n295_), .A2(new_n302_), .A3(KEYINPUT30), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n286_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT31), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n286_), .A3(new_n306_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n309_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n228_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n313_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(new_n227_), .A3(new_n311_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n279_), .A2(new_n280_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n273_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n276_), .A2(KEYINPUT88), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n254_), .A2(new_n257_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n276_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n319_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n323_), .A2(new_n278_), .B1(new_n316_), .B2(new_n314_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n248_), .B1(new_n318_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n268_), .A2(new_n303_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT90), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n289_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n288_), .B(KEYINPUT90), .C1(G183gat), .C2(G190gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n294_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n288_), .A2(new_n301_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT89), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n288_), .A2(new_n301_), .A3(KEYINPUT89), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n300_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n326_), .B1(new_n268_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT20), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT19), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n265_), .B(new_n266_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT95), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n336_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n330_), .A2(KEYINPUT95), .A3(new_n335_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n342_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT20), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT96), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n345_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT95), .B1(new_n330_), .B2(new_n335_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n268_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT96), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT20), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n342_), .A2(new_n303_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n348_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n341_), .B1(new_n355_), .B2(new_n340_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT18), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT98), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n354_), .B(KEYINPUT20), .C1(new_n342_), .C2(new_n336_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n340_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n337_), .A2(KEYINPUT20), .A3(new_n340_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n360_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n356_), .A2(KEYINPUT98), .A3(new_n360_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT27), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n367_), .B(KEYINPUT91), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372_));
  INV_X1    g171(.A(new_n360_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n364_), .A2(new_n365_), .A3(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT92), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n325_), .B1(new_n370_), .B2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n279_), .A2(new_n280_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n317_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n245_), .A2(new_n246_), .B1(new_n366_), .B2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n356_), .A2(new_n380_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(KEYINPUT97), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT97), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n356_), .A2(new_n384_), .A3(new_n380_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n381_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n246_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT93), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n231_), .B(KEYINPUT94), .Z(new_n391_));
  INV_X1    g190(.A(new_n232_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n237_), .A2(new_n392_), .A3(new_n235_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(new_n243_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n246_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n393_), .A2(new_n395_), .B1(new_n396_), .B2(KEYINPUT33), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n390_), .A2(new_n371_), .A3(new_n375_), .A4(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n379_), .B1(new_n386_), .B2(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n377_), .A2(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(KEYINPUT76), .B(G15gat), .Z(new_n401_));
  INV_X1    g200(.A(G22gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G1gat), .A2(G8gat), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n401_), .A2(new_n402_), .B1(KEYINPUT14), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n402_), .B2(new_n401_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G1gat), .B(G8gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT77), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n407_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G29gat), .B(G36gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(G43gat), .B(G50gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n413_), .B(KEYINPUT15), .Z(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n408_), .A2(new_n409_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n413_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G229gat), .A2(G233gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n410_), .A2(new_n413_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n423_), .A2(G229gat), .A3(G233gat), .A4(new_n418_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G113gat), .B(G141gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G169gat), .B(G197gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n428_), .B(KEYINPUT82), .Z(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .A4(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G230gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT7), .ZN(new_n436_));
  INV_X1    g235(.A(G99gat), .ZN(new_n437_));
  INV_X1    g236(.A(G106gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G99gat), .A2(G106gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .A4(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(G85gat), .A2(G92gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(G85gat), .A2(G92gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n445_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT9), .ZN(new_n453_));
  INV_X1    g252(.A(G85gat), .ZN(new_n454_));
  INV_X1    g253(.A(G92gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G85gat), .A2(G92gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n453_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n453_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT64), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT64), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n462_), .B(new_n459_), .C1(new_n448_), .C2(new_n453_), .ZN(new_n463_));
  AND2_X1   g262(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n464_), .A2(new_n465_), .A3(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n442_), .A2(new_n443_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n461_), .A2(new_n463_), .A3(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT66), .B1(new_n452_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n461_), .A2(new_n468_), .A3(new_n463_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT66), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n471_), .B(new_n472_), .C1(new_n451_), .C2(new_n450_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT67), .B(G71gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(G78gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G57gat), .B(G64gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n476_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G78gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n475_), .B(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n479_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n474_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n470_), .A2(new_n485_), .A3(new_n473_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n435_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT68), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n471_), .A2(KEYINPUT69), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n471_), .A2(KEYINPUT69), .ZN(new_n492_));
  INV_X1    g291(.A(new_n452_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT12), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n474_), .A2(new_n486_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n488_), .A2(KEYINPUT70), .A3(new_n495_), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT70), .B1(new_n488_), .B2(new_n495_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n435_), .B(new_n497_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G120gat), .B(G148gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT5), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT71), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G176gat), .B(G204gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n490_), .A2(KEYINPUT72), .A3(new_n500_), .A4(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n487_), .A2(new_n488_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT68), .B1(new_n507_), .B2(new_n435_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n489_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n508_), .A2(new_n500_), .A3(new_n510_), .A4(new_n505_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT72), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n506_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n490_), .A2(new_n500_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n505_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n514_), .A2(KEYINPUT13), .A3(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT73), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(KEYINPUT73), .A3(new_n521_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT37), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n474_), .A2(new_n417_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n494_), .A2(new_n414_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT34), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n528_), .B(new_n529_), .C1(KEYINPUT35), .C2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(KEYINPUT35), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n534_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G190gat), .B(G218gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT74), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT75), .ZN(new_n540_));
  XOR2_X1   g339(.A(G134gat), .B(G162gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(KEYINPUT36), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n542_), .B(KEYINPUT36), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n537_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n527_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT37), .A3(new_n544_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n485_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n410_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G127gat), .B(G155gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT16), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT78), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G183gat), .B(G211gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n559_), .A2(new_n560_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n554_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT80), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n554_), .A2(new_n561_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT79), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n551_), .A2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n400_), .A2(new_n434_), .A3(new_n526_), .A4(new_n568_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n569_), .A2(KEYINPUT99), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(KEYINPUT99), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n248_), .A2(G1gat), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT38), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n400_), .A2(new_n434_), .A3(new_n526_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT100), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n549_), .A2(KEYINPUT100), .A3(new_n544_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(new_n567_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n575_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G1gat), .B1(new_n582_), .B2(new_n248_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n574_), .A2(new_n583_), .ZN(G1324gat));
  AND2_X1   g383(.A1(new_n370_), .A2(new_n376_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(G8gat), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n570_), .A2(new_n571_), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT101), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n575_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(G8gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT39), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT40), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(G1325gat));
  OR3_X1    g394(.A1(new_n569_), .A2(G15gat), .A3(new_n317_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G15gat), .B1(new_n582_), .B2(new_n317_), .ZN(new_n597_));
  XOR2_X1   g396(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n598_));
  AND2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n597_), .A2(new_n598_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n596_), .B1(new_n599_), .B2(new_n600_), .ZN(G1326gat));
  XNOR2_X1  g400(.A(new_n378_), .B(KEYINPUT103), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G22gat), .B1(new_n582_), .B2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT42), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n402_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(new_n569_), .B2(new_n606_), .ZN(G1327gat));
  OAI21_X1  g406(.A(new_n551_), .B1(new_n377_), .B2(new_n399_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT43), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT43), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n610_), .B(new_n551_), .C1(new_n377_), .C2(new_n399_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n525_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT73), .B1(new_n520_), .B2(new_n521_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n567_), .B(new_n434_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT104), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n526_), .A2(new_n617_), .A3(new_n567_), .A4(new_n434_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n612_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n612_), .A2(new_n616_), .A3(KEYINPUT44), .A4(new_n618_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(G29gat), .A3(new_n247_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n567_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n579_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n575_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n248_), .ZN(new_n628_));
  OAI22_X1  g427(.A1(new_n622_), .A2(new_n624_), .B1(G29gat), .B2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT106), .Z(G1328gat));
  OR2_X1    g429(.A1(new_n586_), .A2(G36gat), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT45), .Z(new_n633_));
  NAND3_X1  g432(.A1(new_n621_), .A2(new_n585_), .A3(new_n623_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n634_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT107), .B1(new_n634_), .B2(G36gat), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n633_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT46), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n633_), .B(KEYINPUT46), .C1(new_n635_), .C2(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1329gat));
  INV_X1    g440(.A(new_n317_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n621_), .A2(G43gat), .A3(new_n642_), .A4(new_n623_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n282_), .B1(new_n627_), .B2(new_n317_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(G1330gat));
  INV_X1    g446(.A(new_n627_), .ZN(new_n648_));
  AOI21_X1  g447(.A(G50gat), .B1(new_n648_), .B2(new_n602_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n378_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n623_), .A2(G50gat), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n649_), .B1(new_n651_), .B2(new_n621_), .ZN(G1331gat));
  NOR2_X1   g451(.A1(new_n526_), .A2(new_n434_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n400_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(new_n567_), .A3(new_n551_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n241_), .A3(new_n247_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT109), .ZN(new_n657_));
  INV_X1    g456(.A(new_n581_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n654_), .B2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n653_), .A2(KEYINPUT109), .A3(new_n581_), .A4(new_n400_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(new_n247_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n656_), .B1(new_n662_), .B2(new_n241_), .ZN(G1332gat));
  NOR2_X1   g462(.A1(new_n586_), .A2(G64gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT110), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n655_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n659_), .A2(new_n585_), .A3(new_n660_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT48), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G64gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G64gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT111), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(G1333gat));
  INV_X1    g472(.A(G71gat), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n642_), .A2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT112), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n655_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT49), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n661_), .A2(new_n642_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(G71gat), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT49), .B(new_n674_), .C1(new_n661_), .C2(new_n642_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(G1334gat));
  NAND3_X1  g481(.A1(new_n655_), .A2(new_n482_), .A3(new_n602_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT50), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n661_), .A2(new_n602_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(G78gat), .ZN(new_n686_));
  AOI211_X1 g485(.A(KEYINPUT50), .B(new_n482_), .C1(new_n661_), .C2(new_n602_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(G1335gat));
  NOR3_X1   g487(.A1(new_n654_), .A2(new_n625_), .A3(new_n579_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n454_), .A3(new_n247_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n526_), .A2(new_n625_), .A3(new_n434_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n612_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G85gat), .B1(new_n692_), .B2(new_n248_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(G1336gat));
  NAND3_X1  g493(.A1(new_n689_), .A2(new_n455_), .A3(new_n585_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G92gat), .B1(new_n692_), .B2(new_n586_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1337gat));
  NOR3_X1   g496(.A1(new_n317_), .A2(new_n465_), .A3(new_n464_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n689_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n612_), .A2(new_n642_), .A3(new_n691_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT113), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n700_), .A2(new_n701_), .A3(G99gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n700_), .B2(G99gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT51), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(KEYINPUT114), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n704_), .B(new_n706_), .ZN(G1338gat));
  NAND3_X1  g506(.A1(new_n612_), .A2(new_n650_), .A3(new_n691_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(G106gat), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n709_), .A2(KEYINPUT52), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(KEYINPUT52), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n689_), .A2(new_n438_), .A3(new_n650_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT115), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(new_n713_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n710_), .B(new_n711_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g516(.A1(new_n585_), .A2(new_n248_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n318_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n433_), .B1(new_n506_), .B2(new_n513_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT55), .B(new_n497_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n435_), .A2(KEYINPUT118), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT55), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n500_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n488_), .A2(new_n495_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT70), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n488_), .A2(KEYINPUT70), .A3(new_n495_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n723_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n731_), .A2(KEYINPUT55), .A3(new_n497_), .A4(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n726_), .A3(new_n733_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n734_), .A2(KEYINPUT56), .A3(new_n516_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT56), .B1(new_n734_), .B2(new_n516_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n721_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT119), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT119), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n721_), .B(new_n739_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n423_), .A2(new_n418_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n420_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n419_), .B(KEYINPUT120), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(new_n420_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n428_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n421_), .A2(new_n424_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n746_), .A2(new_n428_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n518_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n738_), .A2(new_n740_), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT57), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n579_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(new_n579_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n745_), .A2(new_n747_), .B1(new_n513_), .B2(new_n506_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT121), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n736_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n734_), .A2(KEYINPUT56), .A3(new_n516_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n736_), .B2(new_n755_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT122), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n551_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n752_), .A2(new_n753_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT123), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n750_), .A2(new_n579_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT57), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n750_), .A2(new_n751_), .A3(new_n579_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n764_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n551_), .A3(new_n762_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(KEYINPUT123), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n625_), .B1(new_n767_), .B2(new_n774_), .ZN(new_n775_));
  XOR2_X1   g574(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n776_));
  NAND4_X1  g575(.A1(new_n520_), .A2(new_n625_), .A3(new_n433_), .A4(new_n521_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT116), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n551_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n777_), .B2(KEYINPUT116), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n776_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n777_), .A2(KEYINPUT116), .ZN(new_n783_));
  INV_X1    g582(.A(new_n776_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n783_), .A2(new_n780_), .A3(new_n778_), .A4(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n720_), .B1(new_n775_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(G113gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n434_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n567_), .B2(new_n765_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n791_), .A2(KEYINPUT59), .A3(new_n719_), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n433_), .B(new_n792_), .C1(new_n787_), .C2(KEYINPUT59), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n790_), .B1(new_n793_), .B2(new_n789_), .ZN(G1340gat));
  NOR2_X1   g593(.A1(new_n613_), .A2(new_n614_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT60), .ZN(new_n796_));
  INV_X1    g595(.A(G120gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n788_), .A2(new_n799_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n526_), .B(new_n792_), .C1(new_n787_), .C2(KEYINPUT59), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n797_), .ZN(G1341gat));
  INV_X1    g601(.A(G127gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n788_), .A2(new_n803_), .A3(new_n625_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n567_), .B(new_n792_), .C1(new_n787_), .C2(KEYINPUT59), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n803_), .ZN(G1342gat));
  INV_X1    g605(.A(G134gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n788_), .A2(new_n807_), .A3(new_n580_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n780_), .B(new_n792_), .C1(new_n787_), .C2(KEYINPUT59), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n807_), .ZN(G1343gat));
  INV_X1    g609(.A(new_n324_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n765_), .A2(new_n766_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT123), .B1(new_n771_), .B2(new_n773_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n567_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n786_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n718_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n203_), .A3(new_n434_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G141gat), .B1(new_n817_), .B2(new_n433_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1344gat));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n204_), .A3(new_n795_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G148gat), .B1(new_n817_), .B2(new_n526_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1345gat));
  XNOR2_X1  g623(.A(KEYINPUT61), .B(G155gat), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n817_), .B2(new_n567_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n816_), .A2(new_n625_), .A3(new_n718_), .A4(new_n825_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1346gat));
  OAI21_X1  g628(.A(G162gat), .B1(new_n817_), .B2(new_n780_), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n579_), .A2(G162gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n817_), .B2(new_n831_), .ZN(G1347gat));
  NOR3_X1   g631(.A1(new_n586_), .A2(new_n247_), .A3(new_n317_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n603_), .ZN(new_n834_));
  NOR4_X1   g633(.A1(new_n791_), .A2(KEYINPUT124), .A3(new_n433_), .A4(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n765_), .A2(new_n567_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n834_), .B1(new_n815_), .B2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n838_), .B2(new_n434_), .ZN(new_n839_));
  OAI21_X1  g638(.A(G169gat), .B1(new_n835_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT62), .B(G169gat), .C1(new_n835_), .C2(new_n839_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n838_), .A2(new_n434_), .A3(new_n292_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n842_), .A2(new_n843_), .A3(new_n844_), .ZN(G1348gat));
  AOI21_X1  g644(.A(new_n650_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n833_), .A2(G176gat), .A3(new_n795_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n838_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n293_), .B1(new_n849_), .B2(new_n526_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(KEYINPUT125), .A3(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1349gat));
  NOR3_X1   g654(.A1(new_n849_), .A2(new_n567_), .A3(new_n296_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n846_), .A2(new_n625_), .A3(new_n833_), .ZN(new_n857_));
  INV_X1    g656(.A(G183gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(G1350gat));
  OAI21_X1  g658(.A(G190gat), .B1(new_n849_), .B2(new_n780_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n838_), .A2(new_n580_), .A3(new_n297_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1351gat));
  NOR2_X1   g661(.A1(new_n586_), .A2(new_n247_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n324_), .B(new_n863_), .C1(new_n775_), .C2(new_n786_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n433_), .ZN(new_n865_));
  INV_X1    g664(.A(G197gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1352gat));
  INV_X1    g666(.A(new_n864_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n526_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n868_), .B(new_n869_), .C1(KEYINPUT126), .C2(G204gat), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n871_));
  INV_X1    g670(.A(G204gat), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n871_), .B(new_n872_), .C1(new_n864_), .C2(new_n526_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n870_), .A2(new_n873_), .ZN(G1353gat));
  NOR2_X1   g673(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n864_), .B2(new_n567_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT63), .B(G211gat), .Z(new_n877_));
  NAND4_X1  g676(.A1(new_n816_), .A2(new_n625_), .A3(new_n863_), .A4(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n876_), .B1(new_n878_), .B2(KEYINPUT127), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT127), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n864_), .A2(new_n567_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n877_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1354gat));
  OAI21_X1  g682(.A(G218gat), .B1(new_n864_), .B2(new_n780_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n579_), .A2(G218gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n864_), .B2(new_n885_), .ZN(G1355gat));
endmodule


