//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  OR2_X1    g002(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n203_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT79), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT23), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n218_));
  AOI21_X1  g017(.A(G176gat), .B1(new_n204_), .B2(new_n205_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(new_n203_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n209_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n202_), .A2(KEYINPUT24), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  MUX2_X1   g027(.A(new_n227_), .B(KEYINPUT24), .S(new_n228_), .Z(new_n229_));
  AND3_X1   g028(.A1(new_n210_), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT78), .B1(new_n210_), .B2(KEYINPUT23), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n213_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT77), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n226_), .A2(new_n229_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n221_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT31), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n235_), .B(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G71gat), .B(G99gat), .Z(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G120gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G113gat), .ZN(new_n242_));
  INV_X1    g041(.A(G113gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G120gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G127gat), .ZN(new_n246_));
  INV_X1    g045(.A(G134gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G127gat), .A2(G134gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n248_), .A2(new_n242_), .A3(new_n244_), .A4(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G15gat), .B(G43gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT80), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n255_), .B(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n240_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n240_), .A2(new_n258_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G155gat), .ZN(new_n263_));
  INV_X1    g062(.A(G162gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT83), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT1), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT83), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(G155gat), .B2(G162gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(G155gat), .A3(G162gat), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n265_), .A2(new_n267_), .A3(new_n269_), .A4(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G141gat), .ZN(new_n273_));
  INV_X1    g072(.A(G148gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT82), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(G141gat), .B2(G148gat), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n272_), .A2(new_n275_), .A3(new_n276_), .A4(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT3), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n276_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n281_), .A2(new_n283_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n265_), .A2(new_n269_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(new_n266_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n279_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G78gat), .B(G106gat), .Z(new_n291_));
  XOR2_X1   g090(.A(new_n290_), .B(new_n291_), .Z(new_n292_));
  INV_X1    g091(.A(G197gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT85), .B1(new_n293_), .B2(G204gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295_));
  INV_X1    g094(.A(G204gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(G197gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(G204gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT86), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n296_), .A2(G197gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT86), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n298_), .A2(new_n300_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G211gat), .ZN(new_n305_));
  INV_X1    g104(.A(G218gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G211gat), .A2(G218gat), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n304_), .A2(KEYINPUT21), .A3(new_n307_), .A4(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n304_), .A2(KEYINPUT21), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT84), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G197gat), .B(G204gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT21), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n293_), .A2(G204gat), .ZN(new_n315_));
  OAI211_X1 g114(.A(KEYINPUT84), .B(KEYINPUT21), .C1(new_n315_), .C2(new_n301_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n307_), .A2(new_n308_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n309_), .B1(new_n310_), .B2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n275_), .A2(new_n278_), .A3(new_n276_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n267_), .A2(new_n271_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n287_), .B2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n265_), .A2(new_n269_), .A3(new_n266_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n284_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n285_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n323_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT29), .B1(new_n322_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n319_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G228gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT28), .ZN(new_n334_));
  XOR2_X1   g133(.A(G22gat), .B(G50gat), .Z(new_n335_));
  XOR2_X1   g134(.A(new_n334_), .B(new_n335_), .Z(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(new_n331_), .A3(new_n319_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n292_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n292_), .B1(new_n339_), .B2(new_n337_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G57gat), .B(G85gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n253_), .B1(new_n322_), .B2(new_n330_), .ZN(new_n351_));
  AND4_X1   g150(.A1(new_n248_), .A2(new_n242_), .A3(new_n244_), .A4(new_n249_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n242_), .A2(new_n244_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n279_), .A2(new_n354_), .A3(new_n288_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(KEYINPUT89), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT89), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n279_), .A2(new_n354_), .A3(new_n357_), .A4(new_n288_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n350_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n351_), .A2(KEYINPUT4), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n358_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(KEYINPUT4), .ZN(new_n362_));
  AOI211_X1 g161(.A(new_n348_), .B(new_n359_), .C1(new_n362_), .C2(new_n350_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT91), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT33), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n232_), .A2(KEYINPUT87), .A3(new_n216_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT87), .B1(new_n232_), .B2(new_n216_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n208_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n307_), .A2(KEYINPUT21), .A3(new_n308_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n299_), .B(new_n302_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n298_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n313_), .A3(new_n298_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n229_), .A2(new_n224_), .A3(new_n214_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n368_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT88), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT88), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n368_), .A2(new_n374_), .A3(new_n378_), .A4(new_n375_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT19), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT20), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n235_), .B2(new_n319_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n377_), .A2(new_n379_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(G92gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT18), .B(G64gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n374_), .B1(new_n368_), .B2(new_n375_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT20), .B1(new_n235_), .B2(new_n319_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n381_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n385_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n385_), .B2(new_n393_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n362_), .A2(new_n349_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT92), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n362_), .A2(KEYINPUT92), .A3(new_n349_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n361_), .A2(new_n350_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n348_), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n361_), .A2(KEYINPUT4), .ZN(new_n403_));
  INV_X1    g202(.A(new_n360_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n350_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n359_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n347_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(KEYINPUT91), .A3(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n365_), .A2(new_n396_), .A3(new_n402_), .A4(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n412_), .A2(new_n349_), .A3(new_n360_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n348_), .B1(new_n413_), .B2(new_n359_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n407_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n391_), .A2(new_n392_), .A3(new_n381_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n235_), .B2(new_n319_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n382_), .B1(new_n419_), .B2(new_n376_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n416_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT93), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n416_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n385_), .A2(new_n393_), .A3(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(KEYINPUT93), .B(new_n416_), .C1(new_n417_), .C2(new_n420_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n415_), .A2(new_n423_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n342_), .B1(new_n410_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n389_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n385_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT27), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT94), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n342_), .A2(new_n414_), .A3(new_n407_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT94), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n429_), .A2(new_n430_), .A3(new_n434_), .A4(KEYINPUT27), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT27), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n437_));
  AND4_X1   g236(.A1(new_n432_), .A2(new_n433_), .A3(new_n435_), .A4(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n262_), .B1(new_n428_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT95), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n437_), .A2(new_n435_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n432_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n415_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n262_), .A2(new_n342_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(KEYINPUT95), .B(new_n262_), .C1(new_n428_), .C2(new_n438_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n441_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT76), .ZN(new_n450_));
  XOR2_X1   g249(.A(G15gat), .B(G22gat), .Z(new_n451_));
  XOR2_X1   g250(.A(KEYINPUT71), .B(G1gat), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G8gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(new_n453_), .B2(KEYINPUT14), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G1gat), .B(G8gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n454_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G29gat), .B(G36gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(G50gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT68), .B(G43gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n457_), .B(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G229gat), .A2(G233gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT74), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n463_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n459_), .A2(new_n460_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n459_), .A2(new_n460_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT15), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT15), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n461_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n471_), .A3(new_n457_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n468_), .B2(new_n457_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n464_), .B1(new_n465_), .B2(new_n473_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n462_), .A2(KEYINPUT74), .A3(new_n463_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n450_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G113gat), .B(G141gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G197gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT75), .B(G169gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n450_), .B(new_n480_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT9), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(G85gat), .A3(G92gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT10), .B(G99gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G85gat), .B(G92gat), .ZN(new_n488_));
  OAI221_X1 g287(.A(new_n486_), .B1(new_n487_), .B2(G106gat), .C1(new_n485_), .C2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n490_));
  AND2_X1   g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n488_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n495_), .B(KEYINPUT7), .Z(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n497_), .A2(KEYINPUT8), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(KEYINPUT8), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n493_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G71gat), .B(G78gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G57gat), .B(G64gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(KEYINPUT11), .B2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(KEYINPUT11), .B2(new_n502_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n501_), .A3(KEYINPUT11), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n507_));
  NOR2_X1   g306(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n508_));
  OAI22_X1  g307(.A1(new_n500_), .A2(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n493_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n497_), .A2(KEYINPUT8), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n497_), .A2(KEYINPUT8), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n506_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n513_), .B(new_n514_), .C1(KEYINPUT66), .C2(KEYINPUT12), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G230gat), .A2(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n500_), .B2(new_n506_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n509_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n510_), .B(new_n506_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT65), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n500_), .A2(new_n506_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n519_), .B1(new_n524_), .B2(new_n516_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G176gat), .B(G204gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(G120gat), .B(G148gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n519_), .B(new_n530_), .C1(new_n524_), .C2(new_n516_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n534_), .A2(KEYINPUT13), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(KEYINPUT13), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n449_), .A2(new_n484_), .A3(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n513_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT34), .ZN(new_n541_));
  OAI22_X1  g340(.A1(new_n513_), .A2(new_n468_), .B1(KEYINPUT35), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n539_), .A2(new_n542_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G134gat), .B(G162gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(KEYINPUT36), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n545_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n550_), .B(KEYINPUT36), .ZN(new_n555_));
  INV_X1    g354(.A(new_n553_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n555_), .B1(new_n556_), .B2(new_n546_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(KEYINPUT70), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(new_n558_), .B2(KEYINPUT37), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n554_), .A2(KEYINPUT69), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT69), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n547_), .A2(new_n565_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n566_), .A3(new_n557_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n561_), .A2(new_n563_), .B1(KEYINPUT37), .B2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G127gat), .B(G155gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(new_n305_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT16), .B(G183gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(KEYINPUT17), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n457_), .B(new_n574_), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(new_n506_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n572_), .A2(KEYINPUT17), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT73), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT72), .ZN(new_n581_));
  AOI211_X1 g380(.A(new_n573_), .B(new_n580_), .C1(new_n581_), .C2(new_n577_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n572_), .B1(new_n581_), .B2(KEYINPUT17), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n576_), .A2(KEYINPUT73), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n568_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n538_), .A2(new_n587_), .ZN(new_n588_));
  OR3_X1    g387(.A1(new_n588_), .A2(new_n452_), .A3(new_n445_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT38), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n586_), .A2(new_n559_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n538_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G1gat), .B1(new_n593_), .B2(new_n445_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n589_), .A2(new_n590_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(new_n594_), .A3(new_n595_), .ZN(G1324gat));
  OR3_X1    g395(.A1(new_n588_), .A2(G8gat), .A3(new_n444_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G8gat), .B1(new_n593_), .B2(new_n444_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n598_), .A2(KEYINPUT39), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(KEYINPUT39), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n597_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g401(.A1(new_n588_), .A2(G15gat), .A3(new_n262_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G15gat), .B1(new_n593_), .B2(new_n262_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT96), .B(KEYINPUT41), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n605_), .A2(new_n606_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n603_), .B1(new_n607_), .B2(new_n608_), .ZN(G1326gat));
  INV_X1    g408(.A(new_n342_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G22gat), .B1(new_n593_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT42), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n610_), .A2(G22gat), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n612_), .B1(new_n588_), .B2(new_n613_), .ZN(G1327gat));
  NOR2_X1   g413(.A1(new_n585_), .A2(new_n558_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n538_), .A2(new_n615_), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n616_), .A2(G29gat), .A3(new_n445_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n537_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n484_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n618_), .A2(new_n619_), .A3(new_n585_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT43), .ZN(new_n621_));
  AOI211_X1 g420(.A(KEYINPUT97), .B(new_n621_), .C1(new_n449_), .C2(new_n568_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n442_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n407_), .A2(KEYINPUT91), .A3(new_n408_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n408_), .B1(new_n407_), .B2(KEYINPUT91), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT92), .B1(new_n362_), .B2(new_n349_), .ZN(new_n627_));
  NOR4_X1   g426(.A1(new_n412_), .A2(new_n398_), .A3(new_n350_), .A4(new_n360_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n401_), .A2(new_n348_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n630_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n415_), .A2(new_n425_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n423_), .A2(new_n426_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n626_), .A2(new_n631_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n623_), .B1(new_n634_), .B2(new_n342_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT95), .B1(new_n635_), .B2(new_n262_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n448_), .A2(new_n447_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n568_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT43), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n620_), .B1(new_n622_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT44), .B(new_n620_), .C1(new_n622_), .C2(new_n640_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n415_), .A3(new_n644_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n645_), .A2(KEYINPUT98), .A3(G29gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT98), .B1(new_n645_), .B2(G29gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n617_), .B1(new_n646_), .B2(new_n647_), .ZN(G1328gat));
  OR2_X1    g447(.A1(new_n443_), .A2(KEYINPUT100), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n443_), .A2(KEYINPUT100), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n616_), .A2(G36gat), .A3(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT45), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n643_), .A2(new_n443_), .A3(new_n644_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT99), .A3(G36gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT99), .B1(new_n654_), .B2(G36gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT46), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(KEYINPUT46), .B(new_n653_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1329gat));
  NAND3_X1  g460(.A1(new_n643_), .A2(new_n261_), .A3(new_n644_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G43gat), .ZN(new_n663_));
  OR3_X1    g462(.A1(new_n616_), .A2(G43gat), .A3(new_n262_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT47), .Z(G1330gat));
  OR3_X1    g465(.A1(new_n616_), .A2(G50gat), .A3(new_n610_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n643_), .A2(new_n342_), .A3(new_n644_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n668_), .A2(KEYINPUT101), .A3(G50gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT101), .B1(new_n668_), .B2(G50gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n667_), .B1(new_n669_), .B2(new_n670_), .ZN(G1331gat));
  NOR2_X1   g470(.A1(new_n537_), .A2(new_n484_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(new_n449_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n592_), .ZN(new_n674_));
  INV_X1    g473(.A(G57gat), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n445_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n587_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT102), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(new_n445_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n676_), .B1(new_n679_), .B2(new_n675_), .ZN(G1332gat));
  OAI21_X1  g479(.A(G64gat), .B1(new_n674_), .B2(new_n651_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT48), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n651_), .A2(G64gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n678_), .B2(new_n683_), .ZN(G1333gat));
  OAI21_X1  g483(.A(G71gat), .B1(new_n674_), .B2(new_n262_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT49), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n262_), .A2(G71gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n678_), .B2(new_n687_), .ZN(G1334gat));
  OAI21_X1  g487(.A(G78gat), .B1(new_n674_), .B2(new_n610_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT103), .B(KEYINPUT50), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n610_), .A2(G78gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n678_), .B2(new_n692_), .ZN(G1335gat));
  NAND2_X1  g492(.A1(new_n673_), .A2(new_n615_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G85gat), .B1(new_n695_), .B2(new_n415_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n622_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n640_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(KEYINPUT104), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n672_), .A2(new_n586_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n622_), .B2(new_n640_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n699_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n415_), .A2(G85gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n696_), .B1(new_n705_), .B2(new_n706_), .ZN(G1336gat));
  INV_X1    g506(.A(G92gat), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n704_), .A2(new_n708_), .A3(new_n651_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n694_), .B2(new_n444_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT105), .ZN(G1337gat));
  OAI21_X1  g511(.A(G99gat), .B1(new_n704_), .B2(new_n262_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n694_), .A2(new_n487_), .A3(new_n262_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(KEYINPUT106), .B2(KEYINPUT51), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(KEYINPUT106), .A2(KEYINPUT51), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n716_), .B(new_n717_), .Z(G1338gat));
  OAI211_X1 g517(.A(new_n342_), .B(new_n701_), .C1(new_n622_), .C2(new_n640_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G106gat), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT108), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(new_n722_), .A3(G106gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n721_), .A2(KEYINPUT52), .A3(new_n723_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n694_), .A2(G106gat), .A3(new_n610_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT107), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT52), .B1(new_n721_), .B2(new_n723_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT53), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n728_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT53), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n726_), .A4(new_n724_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n729_), .A2(new_n732_), .ZN(G1339gat));
  AOI21_X1  g532(.A(new_n484_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n587_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n587_), .A2(new_n734_), .A3(new_n736_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n474_), .A2(new_n475_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n481_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n473_), .A2(KEYINPUT111), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n463_), .B1(new_n473_), .B2(KEYINPUT111), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n742_), .A2(new_n480_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n746_), .A2(new_n747_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n533_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n509_), .A2(new_n515_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n517_), .B1(new_n522_), .B2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n509_), .A2(new_n515_), .A3(new_n518_), .A4(KEYINPUT55), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n519_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n753_), .A3(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n531_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT113), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n750_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT56), .B1(new_n756_), .B2(new_n531_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n758_), .A2(new_n761_), .A3(KEYINPUT113), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT58), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT58), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n760_), .B2(new_n762_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n766_), .A3(new_n568_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n534_), .A2(new_n749_), .A3(new_n748_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n482_), .A2(new_n483_), .A3(new_n533_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n770_), .B1(new_n758_), .B2(new_n761_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(KEYINPUT110), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773_));
  INV_X1    g572(.A(new_n761_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n757_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n775_), .B2(new_n770_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n768_), .B(new_n558_), .C1(new_n772_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n771_), .A2(KEYINPUT110), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n773_), .A3(new_n770_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n769_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n768_), .B1(new_n781_), .B2(new_n558_), .ZN(new_n782_));
  OAI211_X1 g581(.A(KEYINPUT114), .B(new_n767_), .C1(new_n778_), .C2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n586_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n558_), .B1(new_n772_), .B2(new_n776_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n777_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT114), .B1(new_n787_), .B2(new_n767_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n741_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n789_), .A2(new_n415_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n443_), .A2(new_n262_), .A3(new_n342_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n484_), .A3(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n767_), .B1(new_n778_), .B2(new_n782_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n740_), .B1(new_n793_), .B2(new_n586_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(KEYINPUT115), .A2(KEYINPUT59), .ZN(new_n795_));
  AND2_X1   g594(.A1(KEYINPUT115), .A2(KEYINPUT59), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n791_), .B(new_n415_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n794_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n789_), .A2(new_n415_), .A3(new_n791_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(KEYINPUT59), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n619_), .A2(new_n243_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n243_), .A2(new_n792_), .B1(new_n800_), .B2(new_n801_), .ZN(G1340gat));
  OAI21_X1  g601(.A(new_n241_), .B1(new_n537_), .B2(KEYINPUT60), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n241_), .A2(KEYINPUT60), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n790_), .A2(new_n791_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n537_), .B(new_n798_), .C1(new_n799_), .C2(KEYINPUT59), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n241_), .ZN(G1341gat));
  NAND3_X1  g606(.A1(new_n790_), .A2(new_n791_), .A3(new_n585_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n586_), .A2(new_n246_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n246_), .A2(new_n808_), .B1(new_n800_), .B2(new_n809_), .ZN(G1342gat));
  NAND3_X1  g609(.A1(new_n790_), .A2(new_n791_), .A3(new_n559_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n568_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n247_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n247_), .A2(new_n811_), .B1(new_n800_), .B2(new_n813_), .ZN(G1343gat));
  AOI211_X1 g613(.A(new_n261_), .B(new_n610_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n790_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G141gat), .B1(new_n816_), .B2(new_n619_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n790_), .A2(new_n273_), .A3(new_n484_), .A4(new_n815_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1344gat));
  OAI21_X1  g618(.A(G148gat), .B1(new_n816_), .B2(new_n537_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n790_), .A2(new_n274_), .A3(new_n618_), .A4(new_n815_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1345gat));
  NAND4_X1  g621(.A1(new_n789_), .A2(new_n415_), .A3(new_n585_), .A4(new_n815_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT61), .B(G155gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1346gat));
  NAND4_X1  g624(.A1(new_n789_), .A2(new_n415_), .A3(new_n559_), .A4(new_n815_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(KEYINPUT116), .A3(new_n264_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n812_), .A2(new_n264_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n789_), .A2(new_n415_), .A3(new_n815_), .A4(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT116), .B1(new_n826_), .B2(new_n264_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1347gat));
  NOR3_X1   g631(.A1(new_n651_), .A2(new_n262_), .A3(new_n415_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n610_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT118), .B1(new_n794_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836_));
  INV_X1    g635(.A(new_n834_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n585_), .B1(new_n787_), .B2(new_n767_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n836_), .B(new_n837_), .C1(new_n838_), .C2(new_n740_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n484_), .A2(new_n206_), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(KEYINPUT119), .Z(new_n841_));
  NAND3_X1  g640(.A1(new_n835_), .A2(new_n839_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n833_), .A2(new_n484_), .ZN(new_n843_));
  XOR2_X1   g642(.A(new_n843_), .B(KEYINPUT117), .Z(new_n844_));
  NOR3_X1   g643(.A1(new_n794_), .A2(new_n342_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(G169gat), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT62), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n845_), .A2(KEYINPUT62), .A3(new_n846_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n842_), .B1(new_n849_), .B2(new_n850_), .ZN(G1348gat));
  NAND3_X1  g650(.A1(new_n835_), .A2(new_n618_), .A3(new_n839_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n207_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT120), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n855_), .A3(new_n207_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n834_), .A2(new_n207_), .A3(new_n537_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n854_), .A2(new_n856_), .B1(new_n789_), .B2(new_n857_), .ZN(G1349gat));
  NOR2_X1   g657(.A1(new_n586_), .A2(new_n222_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n835_), .A2(new_n839_), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(G183gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n837_), .B1(new_n838_), .B2(new_n740_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n586_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT121), .ZN(G1350gat));
  NAND2_X1  g664(.A1(new_n559_), .A2(new_n223_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT123), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n835_), .A2(new_n839_), .A3(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n835_), .A2(new_n568_), .A3(new_n839_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n869_), .A2(new_n870_), .A3(G190gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n869_), .B2(G190gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n871_), .B2(new_n872_), .ZN(G1351gat));
  NOR4_X1   g672(.A1(new_n651_), .A2(new_n261_), .A3(new_n610_), .A4(new_n415_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n789_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(G197gat), .B1(new_n875_), .B2(new_n484_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n789_), .A2(G197gat), .A3(new_n484_), .A4(new_n874_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n877_), .A2(KEYINPUT124), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(KEYINPUT124), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n876_), .A2(new_n878_), .A3(new_n879_), .ZN(G1352gat));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n618_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n296_), .A2(KEYINPUT125), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1353gat));
  NAND2_X1  g682(.A1(new_n789_), .A2(new_n874_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  AND2_X1   g684(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n884_), .A2(new_n586_), .A3(new_n885_), .A4(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n884_), .B2(new_n586_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT126), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n890_), .B(new_n885_), .C1(new_n884_), .C2(new_n586_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n887_), .B1(new_n889_), .B2(new_n891_), .ZN(G1354gat));
  AOI21_X1  g691(.A(G218gat), .B1(new_n875_), .B2(new_n559_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n884_), .A2(new_n306_), .A3(new_n812_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1355gat));
endmodule


