//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n946_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n964_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G15gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G22gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n208_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G57gat), .B(G64gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n214_));
  XOR2_X1   g013(.A(G71gat), .B(G78gat), .Z(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n214_), .A2(new_n215_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n211_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G127gat), .B(G155gat), .Z(new_n222_));
  XNOR2_X1  g021(.A(G183gat), .B(G211gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT17), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n226_), .A2(KEYINPUT17), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n221_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT65), .B(KEYINPUT6), .Z(new_n232_));
  INV_X1    g031(.A(G99gat), .ZN(new_n233_));
  INV_X1    g032(.A(G106gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT64), .B(G85gat), .ZN(new_n241_));
  INV_X1    g040(.A(G92gat), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n241_), .A2(KEYINPUT9), .A3(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G85gat), .B(G92gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT9), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT10), .B(G99gat), .Z(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n234_), .ZN(new_n247_));
  AND4_X1   g046(.A1(new_n240_), .A2(new_n243_), .A3(new_n245_), .A4(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G99gat), .A2(G106gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT7), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n244_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT8), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n251_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n239_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n238_), .A2(new_n235_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT8), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n244_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n248_), .B1(new_n254_), .B2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G29gat), .B(G36gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G43gat), .B(G50gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT35), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G232gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT34), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n261_), .A2(new_n264_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n260_), .A2(new_n254_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT66), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n260_), .A2(new_n254_), .A3(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n248_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n264_), .B(KEYINPUT15), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n269_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n268_), .A2(new_n265_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G190gat), .B(G218gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G134gat), .B(G162gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(KEYINPUT36), .ZN(new_n283_));
  OAI221_X1 g082(.A(new_n269_), .B1(new_n265_), .B2(new_n268_), .C1(new_n274_), .C2(new_n276_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n279_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT37), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n279_), .A2(new_n284_), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n282_), .B(KEYINPUT36), .Z(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n286_), .B(new_n287_), .C1(new_n288_), .C2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n289_), .B(KEYINPUT69), .Z(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(new_n279_), .B2(new_n284_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT37), .B1(new_n285_), .B2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n231_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT72), .Z(new_n296_));
  NAND4_X1  g095(.A1(new_n240_), .A2(new_n243_), .A3(new_n245_), .A4(new_n247_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n273_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n272_), .B1(new_n260_), .B2(new_n254_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n218_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT12), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n259_), .B1(new_n258_), .B2(new_n244_), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n252_), .A2(KEYINPUT8), .A3(new_n253_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n218_), .B(new_n297_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT12), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n270_), .A2(new_n297_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n301_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n300_), .A2(new_n303_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G230gat), .A2(G233gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n306_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n311_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G120gat), .B(G148gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G176gat), .B(G204gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n312_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n320_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT13), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n324_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n296_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(KEYINPUT1), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT84), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(G155gat), .B2(G162gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(KEYINPUT84), .A3(new_n334_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n334_), .A2(KEYINPUT1), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n338_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n335_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n334_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n344_), .A2(new_n347_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G22gat), .B(G50gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT28), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n361_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G197gat), .B(G204gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n368_));
  OAI211_X1 g167(.A(KEYINPUT21), .B(new_n366_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n367_), .A2(new_n368_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT21), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n366_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(KEYINPUT21), .B2(new_n367_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n369_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n376_));
  AND2_X1   g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n375_), .B2(KEYINPUT85), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  OAI221_X1 g178(.A(new_n375_), .B1(KEYINPUT85), .B2(new_n377_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n365_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n364_), .B1(new_n381_), .B2(KEYINPUT87), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT88), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT88), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n384_), .B(new_n364_), .C1(new_n381_), .C2(KEYINPUT87), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n380_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n365_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(new_n381_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n383_), .A2(new_n385_), .A3(new_n390_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT91), .B(G85gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT0), .B(G57gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G134gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G127gat), .ZN(new_n401_));
  INV_X1    g200(.A(G127gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G134gat), .ZN(new_n403_));
  INV_X1    g202(.A(G120gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(G113gat), .ZN(new_n405_));
  INV_X1    g204(.A(G113gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G120gat), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n401_), .A2(new_n403_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n401_), .A2(new_n403_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(KEYINPUT82), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n412_));
  AND4_X1   g211(.A1(new_n401_), .A2(new_n403_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(new_n408_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n347_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n342_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(new_n341_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n357_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n411_), .B(new_n414_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n419_), .A2(KEYINPUT4), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT90), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n413_), .A2(new_n408_), .ZN(new_n425_));
  NOR4_X1   g224(.A1(new_n417_), .A2(new_n425_), .A3(new_n418_), .A4(KEYINPUT89), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT89), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n409_), .A2(new_n410_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n359_), .B2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n426_), .B1(new_n429_), .B2(new_n419_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n424_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n355_), .A2(new_n358_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n340_), .A2(KEYINPUT84), .A3(new_n334_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT84), .B1(new_n340_), .B2(new_n334_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n342_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n433_), .B(new_n428_), .C1(new_n436_), .C2(new_n415_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n419_), .A2(KEYINPUT89), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n359_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(KEYINPUT90), .A3(KEYINPUT4), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n423_), .B1(new_n432_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n421_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n430_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n399_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT90), .B1(new_n440_), .B2(KEYINPUT4), .ZN(new_n446_));
  AOI211_X1 g245(.A(new_n424_), .B(new_n431_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n422_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n444_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n399_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT27), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G226gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT19), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G169gat), .A2(G176gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT24), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459_));
  MUX2_X1   g258(.A(new_n458_), .B(KEYINPUT24), .S(new_n459_), .Z(new_n460_));
  NAND2_X1  g259(.A1(G183gat), .A2(G190gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT23), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT25), .B(G183gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT26), .B(G190gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n460_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n462_), .B1(G183gat), .B2(G190gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G169gat), .ZN(new_n469_));
  INV_X1    g268(.A(G176gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n457_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n466_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT20), .B1(new_n473_), .B2(new_n375_), .ZN(new_n474_));
  AND2_X1   g273(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n475_));
  NOR2_X1   g274(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n476_));
  OAI21_X1  g275(.A(G169gat), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT79), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT22), .ZN(new_n480_));
  INV_X1    g279(.A(G169gat), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(KEYINPUT77), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT77), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G169gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(G176gat), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(KEYINPUT79), .B(G169gat), .C1(new_n475_), .C2(new_n476_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT80), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n457_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n487_), .B2(new_n457_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n467_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n463_), .A2(KEYINPUT76), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT25), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT76), .B1(new_n493_), .B2(G183gat), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n492_), .A2(new_n494_), .A3(new_n464_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n460_), .A2(new_n462_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(new_n498_), .ZN(new_n499_));
  AOI211_X1 g298(.A(new_n456_), .B(new_n474_), .C1(new_n499_), .C2(new_n375_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G8gat), .B(G36gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT18), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G64gat), .B(G92gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n456_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n375_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n491_), .A2(new_n498_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n473_), .B2(new_n375_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n505_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n500_), .A2(new_n504_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n504_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n456_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n499_), .A2(new_n375_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n474_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n505_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n512_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n454_), .B1(new_n511_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n507_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n474_), .B1(new_n499_), .B2(new_n375_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(new_n505_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n504_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n514_), .A2(new_n517_), .A3(new_n512_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(KEYINPUT27), .A3(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n394_), .A2(new_n453_), .A3(new_n519_), .A4(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n512_), .A2(KEYINPUT32), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(new_n500_), .B2(new_n510_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n520_), .B(new_n529_), .C1(new_n521_), .C2(new_n505_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n445_), .A2(new_n451_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT33), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n399_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n448_), .A2(new_n449_), .A3(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n420_), .A2(new_n443_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n421_), .B1(new_n430_), .B2(KEYINPUT92), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n440_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n450_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n536_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n504_), .B1(new_n500_), .B2(new_n510_), .ZN(new_n542_));
  AND4_X1   g341(.A1(new_n534_), .A2(new_n541_), .A3(new_n524_), .A4(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n451_), .A2(new_n532_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n531_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n526_), .B1(new_n545_), .B2(new_n394_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n487_), .A2(new_n457_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT80), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n487_), .A2(new_n488_), .A3(new_n457_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n468_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n547_), .B1(new_n551_), .B2(new_n497_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n491_), .A2(KEYINPUT30), .A3(new_n498_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G71gat), .B(G99gat), .ZN(new_n554_));
  INV_X1    g353(.A(G43gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G227gat), .A2(G233gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(G15gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n556_), .B(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n552_), .A2(KEYINPUT81), .A3(new_n553_), .A4(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n411_), .A2(new_n414_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT31), .Z(new_n562_));
  INV_X1    g361(.A(KEYINPUT83), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT81), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n551_), .A2(new_n547_), .A3(new_n497_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT30), .B1(new_n491_), .B2(new_n498_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n552_), .A2(KEYINPUT81), .A3(new_n553_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n559_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n562_), .A2(new_n563_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n565_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n574_), .B1(new_n565_), .B2(new_n572_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n452_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT93), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n519_), .A2(new_n525_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n383_), .A2(new_n385_), .A3(new_n390_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n390_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .A4(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n519_), .A2(new_n392_), .A3(new_n393_), .A4(new_n525_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n565_), .A2(new_n572_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n573_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n565_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n588_), .A2(new_n451_), .A3(new_n445_), .A4(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT93), .B1(new_n586_), .B2(new_n590_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n546_), .A2(new_n578_), .B1(new_n585_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n211_), .A2(new_n275_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n209_), .A2(new_n210_), .A3(new_n264_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT73), .ZN(new_n597_));
  INV_X1    g396(.A(new_n594_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n595_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n264_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT73), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n593_), .A2(new_n602_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n597_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G169gat), .B(G197gat), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n605_), .B(new_n606_), .Z(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n604_), .A2(KEYINPUT74), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT74), .B1(new_n604_), .B2(new_n608_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n597_), .A2(new_n601_), .A3(new_n603_), .A4(new_n607_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT75), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n601_), .A2(new_n603_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT75), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n597_), .A4(new_n607_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n611_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n592_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n333_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT94), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT94), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n622_), .A2(new_n204_), .A3(new_n452_), .A4(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n625_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n332_), .A2(new_n618_), .A3(new_n231_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n288_), .A2(new_n290_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(new_n285_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n592_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n453_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n627_), .A3(new_n634_), .ZN(G1324gat));
  OAI21_X1  g434(.A(G8gat), .B1(new_n633_), .B2(new_n581_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT39), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n519_), .A2(new_n525_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n622_), .A2(new_n205_), .A3(new_n640_), .A4(new_n623_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n636_), .A2(new_n637_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(KEYINPUT39), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n639_), .B(new_n641_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(G1325gat));
  OAI21_X1  g445(.A(G15gat), .B1(new_n633_), .B2(new_n578_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT41), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n620_), .A2(G15gat), .A3(new_n578_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1326gat));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n632_), .B2(new_n394_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT42), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n621_), .A2(new_n651_), .A3(new_n394_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1327gat));
  NAND2_X1  g454(.A1(new_n630_), .A2(new_n231_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n332_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n619_), .A2(new_n657_), .ZN(new_n658_));
  OR3_X1    g457(.A1(new_n658_), .A2(G29gat), .A3(new_n453_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n618_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n331_), .A2(new_n660_), .A3(new_n231_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT97), .B(KEYINPUT43), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n291_), .A2(new_n294_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n531_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n511_), .A2(new_n518_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n544_), .A2(new_n670_), .A3(new_n534_), .A4(new_n541_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n394_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n451_), .B(new_n445_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(new_n640_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n578_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n585_), .A2(new_n591_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n668_), .B1(new_n677_), .B2(KEYINPUT98), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT98), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n676_), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n664_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n291_), .A2(new_n294_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n592_), .A2(KEYINPUT43), .A3(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT44), .B(new_n662_), .C1(new_n681_), .C2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n667_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n291_), .A2(new_n294_), .A3(new_n665_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n592_), .B2(new_n679_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n680_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n663_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n683_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n694_), .A2(KEYINPUT100), .A3(KEYINPUT44), .A4(new_n662_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n662_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n686_), .A2(new_n695_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n452_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n699_), .A2(KEYINPUT101), .A3(G29gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT101), .B1(new_n699_), .B2(G29gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n659_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(G36gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n698_), .B2(new_n640_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n658_), .A2(G36gat), .A3(new_n581_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT45), .ZN(new_n707_));
  OR3_X1    g506(.A1(new_n704_), .A2(new_n705_), .A3(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  NAND3_X1  g509(.A1(new_n698_), .A2(G43gat), .A3(new_n577_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n555_), .B1(new_n658_), .B2(new_n578_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(G1330gat));
  INV_X1    g514(.A(G50gat), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n619_), .A2(new_n716_), .A3(new_n394_), .A4(new_n657_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n661_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n394_), .B1(new_n718_), .B2(KEYINPUT44), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n686_), .B2(new_n695_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n716_), .B1(new_n720_), .B2(KEYINPUT103), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n686_), .A2(new_n695_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n584_), .B1(new_n697_), .B2(new_n696_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT103), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT104), .B1(new_n721_), .B2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT100), .B1(new_n718_), .B2(KEYINPUT44), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n585_), .A2(new_n591_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n534_), .A2(new_n541_), .A3(new_n524_), .A4(new_n542_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n442_), .A2(new_n444_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT33), .B1(new_n730_), .B2(new_n450_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n584_), .B1(new_n732_), .B2(new_n531_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n577_), .B1(new_n733_), .B2(new_n526_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT98), .B1(new_n728_), .B2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n680_), .A3(new_n689_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n683_), .B1(new_n736_), .B2(new_n663_), .ZN(new_n737_));
  NOR4_X1   g536(.A1(new_n737_), .A2(new_n685_), .A3(new_n696_), .A4(new_n661_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT103), .B(new_n723_), .C1(new_n727_), .C2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G50gat), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n724_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n717_), .B1(new_n726_), .B2(new_n742_), .ZN(G1331gat));
  NOR4_X1   g542(.A1(new_n296_), .A2(new_n592_), .A3(new_n660_), .A4(new_n331_), .ZN(new_n744_));
  INV_X1    g543(.A(G57gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n452_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n231_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n631_), .A2(new_n618_), .A3(new_n332_), .A4(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n452_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n746_), .B1(new_n751_), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g551(.A(G64gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n744_), .A2(new_n753_), .A3(new_n640_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n750_), .A2(new_n640_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G64gat), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT48), .B(new_n753_), .C1(new_n750_), .C2(new_n640_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT106), .ZN(G1333gat));
  INV_X1    g559(.A(G71gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n750_), .B2(new_n577_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT49), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n744_), .A2(new_n761_), .A3(new_n577_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1334gat));
  INV_X1    g564(.A(G78gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n750_), .B2(new_n394_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n744_), .A2(new_n766_), .A3(new_n394_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1335gat));
  NOR4_X1   g570(.A1(new_n592_), .A2(new_n660_), .A3(new_n331_), .A4(new_n656_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n452_), .ZN(new_n773_));
  NOR4_X1   g572(.A1(new_n737_), .A2(new_n660_), .A3(new_n331_), .A4(new_n747_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n453_), .A2(new_n241_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(G1336gat));
  NAND3_X1  g575(.A1(new_n772_), .A2(new_n242_), .A3(new_n640_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n774_), .A2(new_n640_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n242_), .ZN(G1337gat));
  AOI21_X1  g578(.A(new_n233_), .B1(new_n774_), .B2(new_n577_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n577_), .A2(new_n246_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n772_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT108), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n782_), .A2(new_n783_), .A3(KEYINPUT51), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT51), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n783_), .A2(KEYINPUT51), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n782_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n784_), .A2(new_n787_), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n772_), .A2(new_n234_), .A3(new_n394_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n774_), .A2(new_n394_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(G106gat), .ZN(new_n792_));
  AOI211_X1 g591(.A(KEYINPUT52), .B(new_n234_), .C1(new_n774_), .C2(new_n394_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n789_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  NAND2_X1  g597(.A1(new_n577_), .A2(new_n452_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(new_n586_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802_));
  INV_X1    g601(.A(new_n682_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n613_), .A2(new_n616_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n593_), .A2(new_n595_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n594_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n807_), .B2(new_n806_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n594_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n608_), .A3(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n805_), .A2(new_n321_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n320_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n310_), .A2(KEYINPUT55), .A3(new_n311_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT12), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n261_), .B2(new_n218_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n261_), .A2(new_n218_), .ZN(new_n817_));
  OAI22_X1  g616(.A1(new_n274_), .A2(new_n302_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n314_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n310_), .B2(new_n311_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n814_), .B(new_n819_), .C1(new_n820_), .C2(KEYINPUT111), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n818_), .B2(new_n314_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n813_), .B1(new_n821_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n812_), .B1(new_n826_), .B2(KEYINPUT56), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n820_), .A2(KEYINPUT111), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n824_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n814_), .A4(new_n819_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n813_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n804_), .B1(new_n827_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n803_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n804_), .B(KEYINPUT58), .C1(new_n827_), .C2(new_n832_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n802_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n826_), .A2(KEYINPUT56), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n831_), .B1(new_n830_), .B2(new_n813_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n812_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT58), .B1(new_n840_), .B2(new_n804_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n833_), .A2(new_n834_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(KEYINPUT115), .A4(new_n803_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n321_), .B1(new_n611_), .B2(new_n617_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(KEYINPUT112), .B2(new_n839_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT56), .B1(new_n826_), .B2(KEYINPUT112), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n324_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n805_), .A2(new_n811_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n846_), .A2(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n844_), .B1(new_n851_), .B2(new_n630_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n850_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n826_), .A2(KEYINPUT112), .A3(KEYINPUT56), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n660_), .A2(new_n854_), .A3(new_n321_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n855_), .B2(new_n847_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n630_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(KEYINPUT57), .A3(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n837_), .A2(new_n843_), .A3(new_n852_), .A4(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n231_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n660_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT110), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n295_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n863_), .B2(new_n295_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n862_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n867_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n865_), .A3(new_n861_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n801_), .B1(new_n860_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n801_), .A2(KEYINPUT59), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n851_), .A2(new_n844_), .A3(new_n630_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n856_), .B2(new_n857_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n841_), .A2(new_n803_), .A3(new_n842_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n747_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n868_), .A2(new_n870_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n875_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n874_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G113gat), .B1(new_n883_), .B2(new_n618_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n872_), .A2(new_n406_), .A3(new_n660_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1340gat));
  OAI211_X1 g685(.A(new_n332_), .B(new_n882_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G120gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n404_), .B1(new_n331_), .B2(KEYINPUT60), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n872_), .B(new_n889_), .C1(KEYINPUT60), .C2(new_n404_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT116), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n888_), .A2(new_n893_), .A3(new_n890_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1341gat));
  AOI21_X1  g694(.A(G127gat), .B1(new_n872_), .B2(new_n747_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n883_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n747_), .A2(G127gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT117), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n896_), .B1(new_n897_), .B2(new_n899_), .ZN(G1342gat));
  OAI21_X1  g699(.A(G134gat), .B1(new_n883_), .B2(new_n682_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n872_), .A2(new_n400_), .A3(new_n630_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1343gat));
  AOI21_X1  g702(.A(new_n577_), .B1(new_n860_), .B2(new_n871_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n584_), .A2(new_n640_), .A3(new_n453_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n618_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT118), .B(G141gat), .Z(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1344gat));
  NOR2_X1   g708(.A1(new_n906_), .A2(new_n331_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT119), .B(G148gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1345gat));
  NAND2_X1  g711(.A1(new_n860_), .A2(new_n871_), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n913_), .A2(new_n578_), .A3(new_n905_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(new_n915_), .A3(new_n747_), .ZN(new_n916_));
  OAI21_X1  g715(.A(KEYINPUT120), .B1(new_n906_), .B2(new_n231_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT61), .B(G155gat), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n916_), .A2(new_n917_), .A3(new_n919_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1346gat));
  AND3_X1   g722(.A1(new_n914_), .A2(G162gat), .A3(new_n689_), .ZN(new_n924_));
  AOI21_X1  g723(.A(G162gat), .B1(new_n914_), .B2(new_n630_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1347gat));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n579_), .A2(new_n640_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(KEYINPUT121), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(new_n394_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n930_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n618_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n927_), .B1(new_n932_), .B2(new_n481_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n469_), .ZN(new_n934_));
  OAI211_X1 g733(.A(KEYINPUT62), .B(G169gat), .C1(new_n931_), .C2(new_n618_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n933_), .A2(new_n934_), .A3(new_n935_), .ZN(G1348gat));
  OAI21_X1  g735(.A(new_n470_), .B1(new_n931_), .B2(new_n331_), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n937_), .A2(KEYINPUT122), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(KEYINPUT122), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n394_), .B1(new_n860_), .B2(new_n871_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n929_), .A2(new_n470_), .A3(new_n331_), .ZN(new_n941_));
  AOI22_X1  g740(.A1(new_n938_), .A2(new_n939_), .B1(new_n940_), .B2(new_n941_), .ZN(G1349gat));
  NOR3_X1   g741(.A1(new_n931_), .A2(new_n463_), .A3(new_n231_), .ZN(new_n943_));
  INV_X1    g742(.A(G183gat), .ZN(new_n944_));
  INV_X1    g743(.A(new_n929_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n940_), .A2(new_n747_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n943_), .B1(new_n944_), .B2(new_n946_), .ZN(G1350gat));
  OAI211_X1 g746(.A(new_n803_), .B(new_n930_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n948_), .A2(new_n949_), .A3(G190gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n948_), .B2(G190gat), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n630_), .A2(new_n464_), .ZN(new_n952_));
  OAI22_X1  g751(.A1(new_n950_), .A2(new_n951_), .B1(new_n931_), .B2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  OAI221_X1 g754(.A(KEYINPUT124), .B1(new_n931_), .B2(new_n952_), .C1(new_n950_), .C2(new_n951_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n955_), .A2(new_n956_), .ZN(G1351gat));
  NOR2_X1   g756(.A1(new_n581_), .A2(new_n673_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n904_), .A2(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n660_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g761(.A1(new_n959_), .A2(new_n331_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(KEYINPUT125), .B(G204gat), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1353gat));
  NOR2_X1   g764(.A1(new_n959_), .A2(new_n231_), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n966_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n967_));
  XOR2_X1   g766(.A(KEYINPUT63), .B(G211gat), .Z(new_n968_));
  AOI21_X1  g767(.A(new_n967_), .B1(new_n966_), .B2(new_n968_), .ZN(G1354gat));
  XNOR2_X1  g768(.A(KEYINPUT127), .B(G218gat), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n959_), .A2(new_n682_), .A3(new_n970_), .ZN(new_n971_));
  OR3_X1    g770(.A1(new_n959_), .A2(KEYINPUT126), .A3(new_n857_), .ZN(new_n972_));
  OAI21_X1  g771(.A(KEYINPUT126), .B1(new_n959_), .B2(new_n857_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n971_), .B1(new_n974_), .B2(new_n970_), .ZN(G1355gat));
endmodule


