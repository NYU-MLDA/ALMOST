//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  OR2_X1    g000(.A1(G57gat), .A2(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G57gat), .A2(G64gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G71gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT66), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G71gat), .ZN(new_n208_));
  INV_X1    g007(.A(G78gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n212_));
  OAI211_X1 g011(.A(KEYINPUT11), .B(new_n204_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n206_), .A2(new_n208_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G78gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n202_), .A2(new_n217_), .A3(new_n203_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n214_), .A2(new_n216_), .A3(new_n218_), .A4(new_n210_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT65), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(KEYINPUT65), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n236_), .A2(KEYINPUT65), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n230_), .A2(new_n234_), .A3(new_n238_), .A4(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT10), .B(G99gat), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n227_), .B(new_n228_), .C1(new_n242_), .C2(G106gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT9), .B1(new_n232_), .B2(new_n233_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT9), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n231_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n244_), .A2(KEYINPUT64), .A3(new_n246_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n243_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n220_), .B1(new_n241_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n243_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n244_), .A2(KEYINPUT64), .A3(new_n246_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT64), .B1(new_n244_), .B2(new_n246_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n213_), .A2(new_n219_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n237_), .A4(new_n240_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n252_), .A2(KEYINPUT12), .A3(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n237_), .A3(new_n240_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n220_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G230gat), .A2(G233gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n252_), .A2(new_n258_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n265_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  INV_X1    g067(.A(G204gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT5), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G176gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n267_), .B(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n273_), .A2(KEYINPUT13), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(KEYINPUT13), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n274_), .A2(KEYINPUT67), .A3(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(G29gat), .A2(G36gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G29gat), .A2(G36gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(G43gat), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G29gat), .ZN(new_n284_));
  INV_X1    g083(.A(G36gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G43gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G29gat), .A2(G36gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n283_), .A2(new_n289_), .A3(G50gat), .ZN(new_n290_));
  AOI21_X1  g089(.A(G50gat), .B1(new_n283_), .B2(new_n289_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT69), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G50gat), .ZN(new_n293_));
  NOR3_X1   g092(.A1(new_n281_), .A2(new_n282_), .A3(G43gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n287_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n283_), .A2(new_n289_), .A3(G50gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n292_), .A2(KEYINPUT15), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT15), .B1(new_n292_), .B2(new_n299_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n260_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT70), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n241_), .A2(new_n251_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n290_), .A2(new_n291_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT35), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G232gat), .A2(G233gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n307_), .B(KEYINPUT68), .Z(new_n308_));
  OR2_X1    g107(.A1(new_n308_), .A2(KEYINPUT34), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(KEYINPUT34), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n304_), .A2(new_n305_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n313_), .B(new_n260_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n303_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n309_), .A2(KEYINPUT35), .A3(new_n310_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT71), .B(G190gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G218gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G134gat), .B(G162gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n322_), .A2(KEYINPUT36), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n312_), .A2(new_n302_), .A3(new_n324_), .A4(new_n316_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n292_), .A2(new_n299_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT15), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n292_), .A2(new_n299_), .A3(KEYINPUT15), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n304_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n311_), .A2(new_n306_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n305_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n331_), .B(new_n316_), .C1(new_n260_), .C2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT72), .B1(new_n330_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n325_), .A2(new_n334_), .ZN(new_n335_));
  AND4_X1   g134(.A1(KEYINPUT73), .A2(new_n318_), .A3(new_n323_), .A4(new_n335_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n315_), .A2(new_n317_), .B1(new_n334_), .B2(new_n325_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT73), .B1(new_n337_), .B2(new_n323_), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n322_), .B(KEYINPUT36), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT74), .ZN(new_n340_));
  OAI22_X1  g139(.A1(new_n336_), .A2(new_n338_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT37), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n318_), .A2(new_n335_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n339_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n339_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT75), .B1(new_n337_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n318_), .A2(new_n323_), .A3(new_n335_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n337_), .A2(KEYINPUT73), .A3(new_n323_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n348_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n342_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G15gat), .B(G22gat), .ZN(new_n358_));
  INV_X1    g157(.A(G1gat), .ZN(new_n359_));
  INV_X1    g158(.A(G8gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT14), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G1gat), .B(G8gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G231gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(new_n220_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT78), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G127gat), .B(G155gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G183gat), .B(G211gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT17), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n368_), .B(new_n375_), .Z(new_n376_));
  INV_X1    g175(.A(new_n367_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n374_), .A3(new_n373_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n280_), .A2(new_n357_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT79), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n364_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n332_), .A2(new_n364_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G229gat), .A2(G233gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT80), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n364_), .B(new_n305_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(new_n385_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G113gat), .B(G141gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G197gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT81), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G169gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n387_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G127gat), .B(G134gat), .ZN(new_n400_));
  INV_X1    g199(.A(G113gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G120gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT31), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT25), .B(G183gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT26), .B(G190gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G169gat), .A2(G176gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(KEYINPUT24), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT82), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G183gat), .A2(G190gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT23), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n411_), .A2(KEYINPUT24), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421_));
  OR2_X1    g220(.A1(G183gat), .A2(G190gat), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n417_), .A2(new_n422_), .B1(G169gat), .B2(G176gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT84), .B(G176gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n425_));
  INV_X1    g224(.A(G169gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n425_), .B1(new_n426_), .B2(KEYINPUT22), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT22), .B(G169gat), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n424_), .B(new_n427_), .C1(new_n428_), .C2(new_n425_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n423_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n420_), .A2(new_n421_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n421_), .B1(new_n420_), .B2(new_n430_), .ZN(new_n433_));
  OAI21_X1  g232(.A(G43gat), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(new_n287_), .A3(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G227gat), .A2(G233gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G15gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G71gat), .B(G99gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n438_), .B(new_n439_), .Z(new_n440_));
  NAND3_X1  g239(.A1(new_n434_), .A2(new_n436_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n407_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n434_), .A2(new_n436_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n440_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(KEYINPUT85), .A3(new_n441_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n406_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n442_), .A2(new_n443_), .A3(new_n407_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(new_n405_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G155gat), .A2(G162gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n455_), .A2(KEYINPUT1), .ZN(new_n456_));
  OR2_X1    g255(.A1(G155gat), .A2(G162gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(KEYINPUT1), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G141gat), .A2(G148gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G141gat), .A2(G148gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n455_), .A2(new_n457_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n455_), .A2(KEYINPUT87), .A3(new_n457_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n461_), .B(KEYINPUT3), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n460_), .B(KEYINPUT2), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n463_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G197gat), .B(G204gat), .Z(new_n474_));
  OR3_X1    g273(.A1(new_n474_), .A2(KEYINPUT88), .A3(KEYINPUT21), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT88), .B1(new_n474_), .B2(KEYINPUT21), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(KEYINPUT21), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G211gat), .B(G218gat), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .A4(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n477_), .A2(new_n478_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT89), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n473_), .A2(KEYINPUT29), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT29), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n463_), .A2(new_n485_), .A3(new_n472_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G22gat), .B(G50gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT28), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G78gat), .B(G106gat), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT90), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n486_), .A2(new_n489_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n492_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n484_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n484_), .B1(new_n497_), .B2(new_n495_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT0), .B(G57gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(G85gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(G1gat), .B(G29gat), .Z(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n404_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n473_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n463_), .A2(new_n404_), .A3(new_n472_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G225gat), .A2(G233gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(KEYINPUT4), .A3(new_n508_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n510_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT4), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n473_), .A2(new_n514_), .A3(new_n506_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n505_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(KEYINPUT92), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n511_), .A2(new_n516_), .A3(new_n505_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AND4_X1   g319(.A1(KEYINPUT92), .A2(new_n511_), .A3(new_n516_), .A4(new_n505_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT18), .B(G64gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G92gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G8gat), .B(G36gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(KEYINPUT20), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n420_), .A2(new_n430_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n481_), .A2(new_n479_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n419_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n428_), .A2(new_n424_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n423_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G226gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT19), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n529_), .A2(new_n534_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n420_), .A2(new_n479_), .A3(new_n481_), .A4(new_n430_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(new_n541_), .A3(KEYINPUT20), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(new_n538_), .ZN(new_n543_));
  OAI211_X1 g342(.A(KEYINPUT32), .B(new_n526_), .C1(new_n539_), .C2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n526_), .A2(KEYINPUT32), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n538_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n540_), .A2(new_n541_), .A3(KEYINPUT20), .A4(new_n538_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n545_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n520_), .A2(new_n522_), .A3(new_n544_), .A4(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n526_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n536_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n551_), .B(new_n547_), .C1(new_n552_), .C2(new_n538_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n526_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n509_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n509_), .A2(new_n556_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n513_), .A3(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n512_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n504_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT33), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n519_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n519_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT33), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n555_), .A2(new_n561_), .A3(new_n563_), .A4(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n500_), .B1(new_n550_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT27), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n553_), .A2(new_n568_), .A3(new_n554_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n554_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n551_), .B1(new_n539_), .B2(new_n543_), .ZN(new_n572_));
  OAI211_X1 g371(.A(KEYINPUT93), .B(new_n526_), .C1(new_n546_), .C2(new_n548_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n569_), .B1(new_n574_), .B2(KEYINPUT27), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n564_), .A2(new_n517_), .A3(KEYINPUT92), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n500_), .B1(new_n576_), .B2(new_n521_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n452_), .B1(new_n567_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(KEYINPUT27), .ZN(new_n580_));
  INV_X1    g379(.A(new_n569_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n500_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT85), .B1(new_n447_), .B2(new_n441_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n405_), .B1(new_n450_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n448_), .A2(new_n406_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n584_), .A2(new_n585_), .B1(new_n522_), .B2(new_n520_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n582_), .A2(KEYINPUT94), .A3(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT94), .B1(new_n586_), .B2(new_n582_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n579_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n382_), .A2(new_n399_), .A3(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n381_), .A2(KEYINPUT79), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n520_), .A2(new_n522_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n592_), .A2(G1gat), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n594_), .A2(new_n595_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT38), .ZN(new_n598_));
  OR3_X1    g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n344_), .B1(new_n343_), .B2(new_n339_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n337_), .A2(KEYINPUT75), .A3(new_n346_), .ZN(new_n601_));
  OAI22_X1  g400(.A1(new_n600_), .A2(new_n601_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT97), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n348_), .A2(new_n353_), .A3(KEYINPUT97), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n399_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n280_), .A2(new_n610_), .A3(new_n380_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n613_), .B(new_n589_), .C1(new_n612_), .C2(new_n611_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n593_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n598_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n599_), .A2(new_n615_), .A3(new_n616_), .ZN(G1324gat));
  INV_X1    g416(.A(new_n592_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n360_), .A3(new_n575_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n575_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n621_), .A2(new_n622_), .A3(G8gat), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n621_), .B2(G8gat), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n619_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g425(.A1(new_n592_), .A2(G15gat), .A3(new_n452_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n614_), .A2(new_n452_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(G15gat), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n629_), .A2(KEYINPUT98), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(KEYINPUT98), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n630_), .A2(KEYINPUT41), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT41), .B1(new_n630_), .B2(new_n631_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n627_), .B1(new_n632_), .B2(new_n633_), .ZN(G1326gat));
  INV_X1    g433(.A(new_n500_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G22gat), .B1(new_n614_), .B2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT99), .B(KEYINPUT42), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT100), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n636_), .B(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n635_), .A2(G22gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT101), .Z(new_n641_));
  OAI21_X1  g440(.A(new_n639_), .B1(new_n592_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1327gat));
  NOR2_X1   g443(.A1(new_n608_), .A2(new_n379_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n280_), .A2(new_n610_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n589_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n593_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n589_), .A2(new_n651_), .A3(new_n357_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n356_), .B(KEYINPUT103), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n589_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n652_), .B1(new_n654_), .B2(new_n651_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n646_), .A3(new_n380_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n284_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n656_), .A2(new_n657_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n593_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n650_), .B1(new_n659_), .B2(new_n661_), .ZN(G1328gat));
  NOR3_X1   g461(.A1(new_n647_), .A2(G36gat), .A3(new_n620_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n658_), .A2(new_n660_), .A3(new_n620_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n285_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT46), .B(new_n665_), .C1(new_n666_), .C2(new_n285_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1329gat));
  OR2_X1    g470(.A1(new_n656_), .A2(new_n657_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n452_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n656_), .A2(new_n657_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n672_), .A2(G43gat), .A3(new_n673_), .A4(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n287_), .B1(new_n647_), .B2(new_n452_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n648_), .B2(new_n500_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n658_), .A2(new_n293_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n660_), .A2(new_n635_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(G1331gat));
  INV_X1    g481(.A(new_n280_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n399_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(new_n589_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n357_), .A2(new_n380_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G57gat), .B1(new_n688_), .B2(new_n649_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n379_), .A3(new_n608_), .ZN(new_n690_));
  INV_X1    g489(.A(G57gat), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n593_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n689_), .A2(new_n692_), .ZN(G1332gat));
  OAI21_X1  g492(.A(G64gat), .B1(new_n690_), .B2(new_n620_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT48), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n620_), .A2(G64gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n687_), .B2(new_n696_), .ZN(G1333gat));
  OAI21_X1  g496(.A(G71gat), .B1(new_n690_), .B2(new_n452_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT49), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n688_), .A2(new_n205_), .A3(new_n673_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1334gat));
  OAI21_X1  g500(.A(G78gat), .B1(new_n690_), .B2(new_n635_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT50), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n688_), .A2(new_n209_), .A3(new_n500_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1335gat));
  NAND2_X1  g504(.A1(new_n685_), .A2(new_n645_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G85gat), .B1(new_n707_), .B2(new_n649_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n589_), .A2(new_n651_), .A3(new_n357_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n651_), .B1(new_n589_), .B2(new_n653_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n380_), .B(new_n684_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(G85gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n708_), .B1(new_n713_), .B2(new_n649_), .ZN(G1336gat));
  AOI21_X1  g513(.A(G92gat), .B1(new_n707_), .B2(new_n575_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n575_), .A2(G92gat), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT105), .Z(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n712_), .B2(new_n717_), .ZN(G1337gat));
  AOI21_X1  g517(.A(new_n222_), .B1(new_n712_), .B2(new_n673_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n706_), .A2(new_n242_), .A3(new_n452_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g521(.A(KEYINPUT53), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n724_));
  OAI21_X1  g523(.A(G106gat), .B1(new_n711_), .B2(new_n635_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT52), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(G106gat), .C1(new_n711_), .C2(new_n635_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n706_), .A2(G106gat), .A3(new_n635_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n724_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT106), .B(new_n730_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n723_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n728_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n655_), .A2(new_n380_), .A3(new_n500_), .A4(new_n684_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n727_), .B1(new_n736_), .B2(G106gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n731_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT106), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n729_), .A2(new_n724_), .A3(new_n731_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(KEYINPUT53), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n734_), .A2(new_n741_), .ZN(G1339gat));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n267_), .A2(new_n272_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n264_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n259_), .A2(new_n745_), .A3(new_n262_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n748_));
  AOI211_X1 g547(.A(KEYINPUT55), .B(new_n745_), .C1(new_n259_), .C2(new_n262_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n750_), .A2(KEYINPUT56), .A3(new_n272_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT56), .B1(new_n750_), .B2(new_n272_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n399_), .B(new_n744_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n386_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n383_), .A2(new_n384_), .A3(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n396_), .B(new_n755_), .C1(new_n388_), .C2(new_n754_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n273_), .A2(new_n398_), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n753_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT57), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT57), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n758_), .A2(new_n604_), .A3(new_n761_), .A4(new_n606_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  INV_X1    g563(.A(new_n746_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n265_), .A2(KEYINPUT55), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n263_), .A2(new_n747_), .A3(new_n264_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n272_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n750_), .A2(KEYINPUT56), .A3(new_n272_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT108), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n750_), .A2(new_n775_), .A3(KEYINPUT56), .A4(new_n272_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n752_), .A2(KEYINPUT109), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n772_), .A2(new_n774_), .A3(new_n776_), .A4(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n744_), .A2(new_n398_), .A3(new_n756_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(KEYINPUT110), .A2(KEYINPUT58), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n778_), .B(new_n779_), .C1(KEYINPUT110), .C2(KEYINPUT58), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n357_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n763_), .A2(KEYINPUT111), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT111), .B1(new_n763_), .B2(new_n784_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(new_n379_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n379_), .A2(new_n610_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(new_n276_), .A3(new_n356_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT54), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n743_), .B1(new_n787_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n763_), .A2(new_n784_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n763_), .A2(KEYINPUT111), .A3(new_n784_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n380_), .A3(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT112), .A3(new_n792_), .ZN(new_n800_));
  NOR4_X1   g599(.A1(new_n452_), .A2(new_n575_), .A3(new_n593_), .A4(new_n500_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT59), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n795_), .A2(new_n380_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n792_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n801_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n399_), .A2(G113gat), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT114), .Z(new_n810_));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n802_), .B(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n399_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n811_), .B1(new_n814_), .B2(new_n401_), .ZN(G1340gat));
  NAND3_X1  g614(.A1(new_n803_), .A2(new_n280_), .A3(new_n807_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n803_), .A2(KEYINPUT116), .A3(new_n280_), .A4(new_n807_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(G120gat), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n403_), .B1(new_n683_), .B2(KEYINPUT60), .ZN(new_n821_));
  XOR2_X1   g620(.A(new_n821_), .B(KEYINPUT115), .Z(new_n822_));
  OAI211_X1 g621(.A(new_n813_), .B(new_n822_), .C1(KEYINPUT60), .C2(new_n403_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1341gat));
  AOI21_X1  g623(.A(G127gat), .B1(new_n813_), .B2(new_n379_), .ZN(new_n825_));
  INV_X1    g624(.A(G127gat), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n808_), .A2(new_n826_), .A3(new_n380_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1342gat));
  AOI21_X1  g627(.A(G134gat), .B1(new_n813_), .B2(new_n609_), .ZN(new_n829_));
  INV_X1    g628(.A(G134gat), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n808_), .A2(new_n830_), .A3(new_n356_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1343gat));
  AND3_X1   g631(.A1(new_n799_), .A2(KEYINPUT112), .A3(new_n792_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT112), .B1(new_n799_), .B2(new_n792_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n620_), .A2(new_n649_), .A3(new_n452_), .A4(new_n500_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT117), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n399_), .A3(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g638(.A1(new_n835_), .A2(new_n280_), .A3(new_n837_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g640(.A(KEYINPUT61), .B(G155gat), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n835_), .A2(new_n379_), .A3(new_n837_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n844_), .A2(new_n845_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n843_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n844_), .A2(new_n845_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n842_), .A3(new_n846_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1346gat));
  NAND4_X1  g651(.A1(new_n835_), .A2(G162gat), .A3(new_n653_), .A4(new_n837_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n794_), .A2(new_n609_), .A3(new_n800_), .A4(new_n837_), .ZN(new_n854_));
  INV_X1    g653(.A(G162gat), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n854_), .A2(KEYINPUT120), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT120), .B1(new_n854_), .B2(new_n855_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n853_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT121), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n860_), .B(new_n853_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1347gat));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n586_), .A2(new_n575_), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n864_), .B(KEYINPUT122), .Z(new_n865_));
  NAND3_X1  g664(.A1(new_n805_), .A2(new_n635_), .A3(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n610_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n426_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n863_), .B1(new_n868_), .B2(KEYINPUT123), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(KEYINPUT123), .B2(new_n868_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n867_), .A2(new_n428_), .ZN(new_n871_));
  OR3_X1    g670(.A1(new_n868_), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(G1348gat));
  NOR3_X1   g672(.A1(new_n833_), .A2(new_n834_), .A3(new_n500_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n865_), .A2(G176gat), .A3(new_n280_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n866_), .A2(new_n683_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n874_), .A2(new_n875_), .B1(new_n876_), .B2(new_n424_), .ZN(G1349gat));
  NOR3_X1   g676(.A1(new_n866_), .A2(new_n380_), .A3(new_n408_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n874_), .A2(new_n379_), .A3(new_n865_), .ZN(new_n879_));
  INV_X1    g678(.A(G183gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(G1350gat));
  OAI21_X1  g680(.A(G190gat), .B1(new_n866_), .B2(new_n356_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n609_), .A2(new_n409_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n866_), .B2(new_n883_), .ZN(G1351gat));
  INV_X1    g683(.A(new_n577_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n673_), .A2(new_n620_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n794_), .A2(new_n885_), .A3(new_n800_), .A4(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n610_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G197gat), .B1(new_n888_), .B2(KEYINPUT124), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n888_), .B2(KEYINPUT124), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892_));
  NOR4_X1   g691(.A1(new_n887_), .A2(new_n892_), .A3(KEYINPUT125), .A4(new_n610_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n889_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(G197gat), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n835_), .A2(new_n399_), .A3(new_n885_), .A4(new_n886_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n892_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n886_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n833_), .A2(new_n834_), .A3(new_n898_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n899_), .A2(KEYINPUT124), .A3(new_n399_), .A4(new_n885_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT125), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n888_), .A2(KEYINPUT124), .A3(new_n890_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n897_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n894_), .A2(new_n903_), .ZN(G1352gat));
  NOR2_X1   g703(.A1(new_n887_), .A2(new_n683_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n269_), .ZN(G1353gat));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n907_));
  INV_X1    g706(.A(G211gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n379_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n887_), .A2(KEYINPUT126), .A3(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT126), .B1(new_n887_), .B2(new_n909_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n907_), .A2(new_n908_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n910_), .A2(new_n907_), .A3(new_n908_), .A4(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1354gat));
  NAND4_X1  g715(.A1(new_n899_), .A2(G218gat), .A3(new_n885_), .A4(new_n357_), .ZN(new_n917_));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n887_), .B2(new_n608_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT127), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n917_), .A2(new_n922_), .A3(new_n919_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1355gat));
endmodule


