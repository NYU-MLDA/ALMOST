//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT36), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT75), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G29gat), .B(G36gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(new_n208_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT6), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT6), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n223_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n222_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n217_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n219_), .A2(new_n221_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n229_), .A2(new_n235_), .A3(new_n231_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT8), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n234_), .A2(KEYINPUT8), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT9), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT9), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT65), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n240_), .B(new_n242_), .C1(G85gat), .C2(G92gat), .ZN(new_n243_));
  OR2_X1    g042(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(G85gat), .A3(new_n245_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n243_), .A2(new_n246_), .B1(KEYINPUT9), .B2(new_n215_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n235_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT10), .B(G99gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT64), .B(G106gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n247_), .A2(new_n248_), .A3(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT69), .B1(new_n238_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n243_), .A2(new_n246_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n251_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n235_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT8), .ZN(new_n260_));
  INV_X1    g059(.A(new_n233_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n261_), .A2(new_n229_), .A3(new_n231_), .A4(new_n223_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n262_), .B2(new_n217_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n236_), .A2(new_n237_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n254_), .B(new_n259_), .C1(new_n263_), .C2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n214_), .B1(new_n253_), .B2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n268_));
  XNOR2_X1  g067(.A(new_n214_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n259_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n248_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(KEYINPUT70), .A3(new_n258_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n234_), .A2(KEYINPUT8), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n264_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n269_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n267_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G232gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n281_), .A2(KEYINPUT35), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT35), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n214_), .B(new_n268_), .Z(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT70), .B1(new_n272_), .B2(new_n258_), .ZN(new_n285_));
  NOR4_X1   g084(.A1(new_n247_), .A2(new_n270_), .A3(new_n251_), .A4(new_n248_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n284_), .B1(new_n287_), .B2(new_n238_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n283_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n278_), .A2(new_n282_), .B1(new_n290_), .B2(new_n281_), .ZN(new_n291_));
  OAI211_X1 g090(.A(KEYINPUT35), .B(new_n281_), .C1(new_n277_), .C2(KEYINPUT74), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n292_), .A2(new_n277_), .A3(new_n267_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n207_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT37), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n254_), .B1(new_n276_), .B2(new_n259_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n238_), .A2(KEYINPUT69), .A3(new_n252_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n288_), .B(new_n282_), .C1(new_n298_), .C2(new_n214_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n292_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n204_), .B(KEYINPUT36), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n278_), .A2(new_n281_), .A3(new_n290_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n294_), .A2(new_n295_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n301_), .A2(new_n305_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n300_), .A2(new_n302_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n295_), .B1(new_n294_), .B2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT77), .B1(new_n304_), .B2(new_n309_), .ZN(new_n310_));
  AND4_X1   g109(.A1(new_n300_), .A2(new_n302_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n207_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT37), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n294_), .A2(new_n295_), .A3(new_n303_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n310_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n320_));
  OR4_X1    g119(.A1(new_n320_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n321_));
  INV_X1    g120(.A(G141gat), .ZN(new_n322_));
  INV_X1    g121(.A(G148gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n320_), .B1(new_n324_), .B2(KEYINPUT3), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT88), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(KEYINPUT3), .B2(new_n324_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(KEYINPUT88), .A3(new_n328_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n326_), .A2(new_n330_), .A3(new_n331_), .A4(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(G155gat), .B2(G162gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n324_), .A2(KEYINPUT85), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n324_), .A2(KEYINPUT85), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT1), .ZN(new_n343_));
  OAI221_X1 g142(.A(new_n327_), .B1(new_n340_), .B2(new_n341_), .C1(new_n336_), .C2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n338_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT29), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT89), .B(G204gat), .ZN(new_n348_));
  OAI211_X1 g147(.A(KEYINPUT21), .B(new_n347_), .C1(new_n348_), .C2(G197gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT21), .ZN(new_n350_));
  INV_X1    g149(.A(G197gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G204gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n350_), .B(new_n352_), .C1(new_n348_), .C2(new_n351_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G211gat), .B(G218gat), .Z(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n349_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT90), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n349_), .A2(new_n353_), .A3(KEYINPUT90), .A4(new_n355_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n352_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(KEYINPUT21), .A3(new_n354_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n346_), .A2(new_n363_), .ZN(new_n364_));
  AND3_X1   g163(.A1(KEYINPUT91), .A2(G228gat), .A3(G233gat), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT91), .B1(G228gat), .B2(G233gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n366_), .B1(new_n364_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n345_), .A2(KEYINPUT29), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT28), .B(G22gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n345_), .A2(KEYINPUT29), .A3(new_n373_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G78gat), .B(G106gat), .ZN(new_n378_));
  INV_X1    g177(.A(G50gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n371_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n370_), .A2(new_n383_), .A3(new_n382_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G92gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT18), .B(G64gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT32), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT20), .ZN(new_n395_));
  INV_X1    g194(.A(new_n362_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n397_));
  INV_X1    g196(.A(G169gat), .ZN(new_n398_));
  INV_X1    g197(.A(G176gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT82), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(G183gat), .A3(G190gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n404_), .A3(KEYINPUT23), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT23), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(G183gat), .ZN(new_n408_));
  INV_X1    g207(.A(G190gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n400_), .B1(new_n411_), .B2(KEYINPUT83), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n405_), .A2(new_n413_), .A3(new_n407_), .A4(new_n410_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT22), .B(G169gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n399_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT24), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(G169gat), .B2(G176gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G169gat), .A2(G176gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT81), .ZN(new_n422_));
  AOI211_X1 g221(.A(new_n418_), .B(new_n400_), .C1(new_n420_), .C2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT26), .B(G190gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT25), .B(G183gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n420_), .A3(new_n418_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n423_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n401_), .A2(new_n406_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n402_), .A2(new_n404_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n431_), .B2(new_n406_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n412_), .A2(new_n417_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n395_), .B1(new_n397_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n406_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n430_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n410_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT94), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n400_), .B(KEYINPUT93), .Z(new_n439_));
  INV_X1    g238(.A(KEYINPUT94), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n432_), .A2(new_n440_), .A3(new_n410_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n438_), .A2(new_n416_), .A3(new_n439_), .A4(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n423_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT92), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n425_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n425_), .A2(new_n444_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n424_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n405_), .A2(new_n407_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n421_), .A2(new_n418_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n443_), .A2(new_n447_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n442_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n363_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G226gat), .A2(G233gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT19), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n434_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT99), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n434_), .A2(new_n452_), .A3(KEYINPUT99), .A4(new_n455_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n451_), .A2(KEYINPUT98), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT98), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n442_), .A2(new_n450_), .A3(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n397_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n417_), .A2(new_n412_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n429_), .A2(new_n432_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n395_), .B1(new_n363_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n455_), .B1(new_n464_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n394_), .B1(new_n460_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G127gat), .B(G134gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G113gat), .B(G120gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n345_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n338_), .A2(new_n473_), .A3(new_n344_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(KEYINPUT4), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G225gat), .A2(G233gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n478_), .B(KEYINPUT95), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT96), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n345_), .A2(new_n481_), .A3(new_n474_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(new_n480_), .A3(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n479_), .A3(new_n476_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(G85gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT0), .B(G57gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n483_), .A2(new_n484_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n434_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n397_), .A2(new_n450_), .A3(new_n442_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n454_), .B1(new_n468_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n393_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n470_), .A2(new_n493_), .A3(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n475_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT97), .B1(new_n501_), .B2(new_n491_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n477_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT97), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n504_), .A3(new_n489_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n392_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n363_), .A2(new_n451_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT20), .B1(new_n397_), .B2(new_n433_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n455_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n392_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n494_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n506_), .A2(new_n507_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT33), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n492_), .A2(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n483_), .A2(KEYINPUT33), .A3(new_n484_), .A4(new_n491_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n388_), .B1(new_n499_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n511_), .B1(new_n460_), .B2(new_n469_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(KEYINPUT27), .A3(new_n507_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n507_), .A2(new_n512_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT27), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT100), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT100), .ZN(new_n525_));
  AOI211_X1 g324(.A(new_n525_), .B(KEYINPUT27), .C1(new_n507_), .C2(new_n512_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n387_), .B(new_n521_), .C1(new_n524_), .C2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n519_), .B1(new_n527_), .B2(new_n493_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT30), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n433_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G15gat), .B(G43gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G227gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n531_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G71gat), .B(G99gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n473_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n535_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n528_), .A2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n510_), .A2(new_n511_), .A3(new_n494_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n511_), .B1(new_n510_), .B2(new_n494_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n523_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n525_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n522_), .A2(KEYINPUT100), .A3(new_n523_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n521_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n538_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n493_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n388_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n319_), .B1(new_n539_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G57gat), .B(G64gat), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n556_), .A2(KEYINPUT11), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(KEYINPUT11), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G71gat), .B(G78gat), .ZN(new_n559_));
  OR3_X1    g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n559_), .A3(KEYINPUT11), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n253_), .A2(new_n266_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n555_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT12), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(KEYINPUT12), .B(new_n564_), .C1(new_n287_), .C2(new_n238_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n568_), .A2(new_n555_), .A3(new_n563_), .A4(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT71), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n564_), .B1(new_n253_), .B2(new_n266_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n567_), .B2(new_n565_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n574_), .A2(KEYINPUT71), .A3(new_n555_), .A4(new_n569_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n566_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G204gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT5), .B(G176gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  AOI211_X1 g381(.A(new_n566_), .B(new_n580_), .C1(new_n572_), .C2(new_n575_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n554_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n566_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n570_), .A2(new_n571_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n570_), .A2(new_n571_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n580_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n576_), .A2(new_n581_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(KEYINPUT13), .A3(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n584_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(G211gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT16), .B(G183gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n594_), .B(new_n595_), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT17), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT79), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G15gat), .B(G22gat), .ZN(new_n599_));
  INV_X1    g398(.A(G1gat), .ZN(new_n600_));
  INV_X1    g399(.A(G8gat), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT14), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G1gat), .B(G8gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT78), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n605_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(new_n564_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n598_), .A2(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT80), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT17), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n609_), .A2(new_n612_), .A3(new_n596_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(KEYINPUT80), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n605_), .B(new_n214_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n605_), .A2(new_n214_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n284_), .B2(new_n605_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620_));
  MUX2_X1   g419(.A(new_n617_), .B(new_n619_), .S(new_n620_), .Z(new_n621_));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G169gat), .B(G197gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n621_), .B(new_n624_), .Z(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n592_), .A2(new_n616_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n553_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n600_), .A3(new_n493_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT38), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n539_), .A2(new_n552_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n291_), .A2(new_n293_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n313_), .B1(new_n301_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT101), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n628_), .A2(new_n632_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G1gat), .B1(new_n637_), .B2(new_n549_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n631_), .A2(new_n638_), .ZN(G1324gat));
  NAND3_X1  g438(.A1(new_n629_), .A2(new_n601_), .A3(new_n546_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n546_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G8gat), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n642_), .A2(KEYINPUT39), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(KEYINPUT39), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(G1325gat));
  INV_X1    g446(.A(G15gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n629_), .A2(new_n648_), .A3(new_n548_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n636_), .B2(new_n548_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n651_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n649_), .B1(new_n655_), .B2(new_n656_), .ZN(G1326gat));
  INV_X1    g456(.A(G22gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n387_), .B(KEYINPUT103), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n636_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT42), .Z(new_n661_));
  NAND3_X1  g460(.A1(new_n629_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1327gat));
  INV_X1    g462(.A(new_n634_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n539_), .B2(new_n552_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n592_), .A2(new_n615_), .A3(new_n626_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n493_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  AOI211_X1 g469(.A(KEYINPUT43), .B(new_n318_), .C1(new_n539_), .C2(new_n552_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n539_), .A2(KEYINPUT104), .A3(new_n552_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n310_), .A2(KEYINPUT105), .A3(new_n317_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT105), .B1(new_n310_), .B2(new_n317_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n545_), .A2(new_n549_), .A3(new_n387_), .A4(new_n521_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n548_), .B1(new_n677_), .B2(new_n519_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n546_), .A2(new_n550_), .A3(new_n387_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n672_), .A2(new_n675_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n671_), .B1(new_n681_), .B2(KEYINPUT43), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n670_), .B1(new_n682_), .B2(new_n666_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n683_), .A2(G29gat), .A3(new_n493_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(new_n671_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(KEYINPUT44), .A3(new_n667_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n669_), .B1(new_n684_), .B2(new_n688_), .ZN(G1328gat));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT106), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT107), .Z(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n668_), .A2(new_n694_), .A3(new_n546_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n668_), .A2(KEYINPUT45), .A3(new_n694_), .A4(new_n546_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n688_), .A2(new_n683_), .A3(new_n546_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(G36gat), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n690_), .A2(KEYINPUT106), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n693_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n702_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n666_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n547_), .B1(new_n705_), .B2(KEYINPUT44), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n694_), .B1(new_n706_), .B2(new_n683_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n692_), .B(new_n704_), .C1(new_n707_), .C2(new_n699_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n703_), .A2(new_n708_), .ZN(G1329gat));
  NAND4_X1  g508(.A1(new_n688_), .A2(new_n683_), .A3(G43gat), .A4(new_n548_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n668_), .A2(new_n548_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n711_), .A2(G43gat), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(G1330gat));
  AOI21_X1  g514(.A(G50gat), .B1(new_n668_), .B2(new_n659_), .ZN(new_n716_));
  AOI211_X1 g515(.A(new_n379_), .B(new_n388_), .C1(new_n705_), .C2(KEYINPUT44), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n683_), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n592_), .A2(new_n626_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n553_), .A2(new_n616_), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G57gat), .B1(new_n720_), .B2(new_n493_), .ZN(new_n721_));
  AND4_X1   g520(.A1(new_n632_), .A2(new_n635_), .A3(new_n719_), .A4(new_n616_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n493_), .A2(G57gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n720_), .A2(new_n725_), .A3(new_n546_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n722_), .B2(new_n546_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT109), .Z(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(KEYINPUT48), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(KEYINPUT48), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(G1333gat));
  INV_X1    g530(.A(G71gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n720_), .A2(new_n732_), .A3(new_n548_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n722_), .B2(new_n548_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT110), .Z(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT49), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(KEYINPUT49), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1334gat));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n722_), .B2(new_n659_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT50), .Z(new_n741_));
  NAND2_X1  g540(.A1(new_n659_), .A2(new_n739_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT111), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n720_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n744_), .ZN(G1335gat));
  NAND2_X1  g544(.A1(new_n584_), .A2(new_n591_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n615_), .A3(new_n625_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n665_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n665_), .A2(KEYINPUT112), .A3(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G85gat), .B1(new_n753_), .B2(new_n493_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n747_), .B(KEYINPUT113), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n682_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n493_), .A2(G85gat), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT114), .Z(new_n759_));
  AOI21_X1  g558(.A(new_n754_), .B1(new_n757_), .B2(new_n759_), .ZN(G1336gat));
  AOI21_X1  g559(.A(G92gat), .B1(new_n753_), .B2(new_n546_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n546_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n757_), .B2(new_n762_), .ZN(G1337gat));
  AOI21_X1  g562(.A(new_n224_), .B1(new_n757_), .B2(new_n548_), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n538_), .B(new_n249_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n766_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n767_), .B(new_n768_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1338gat));
  XNOR2_X1  g572(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n682_), .A2(new_n388_), .A3(new_n756_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT52), .B1(new_n775_), .B2(new_n225_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n687_), .A2(new_n387_), .A3(new_n755_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(G106gat), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n388_), .B(new_n250_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n774_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n774_), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n784_), .B(new_n781_), .C1(new_n776_), .C2(new_n779_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n592_), .A2(new_n616_), .A3(new_n318_), .A4(new_n625_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(KEYINPUT54), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n584_), .A2(new_n591_), .A3(new_n616_), .A4(new_n625_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n319_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(KEYINPUT117), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT54), .B1(new_n319_), .B2(new_n790_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n788_), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT119), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(new_n572_), .B2(new_n575_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n574_), .A2(KEYINPUT55), .A3(new_n555_), .A4(new_n569_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n574_), .A2(new_n569_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n555_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n580_), .B(new_n802_), .C1(new_n803_), .C2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n570_), .A2(new_n808_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n555_), .B1(new_n574_), .B2(new_n569_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n581_), .B1(new_n809_), .B2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n801_), .B1(new_n576_), .B2(new_n581_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n626_), .B(new_n807_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n617_), .A2(new_n620_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n619_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n620_), .ZN(new_n818_));
  MUX2_X1   g617(.A(new_n621_), .B(new_n818_), .S(new_n624_), .Z(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n664_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(KEYINPUT57), .A3(new_n664_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n590_), .B1(new_n813_), .B2(new_n800_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n580_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n819_), .B1(new_n828_), .B2(KEYINPUT56), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n826_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n583_), .B1(new_n828_), .B2(KEYINPUT56), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n813_), .A2(new_n800_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(KEYINPUT58), .A4(new_n819_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(new_n319_), .A3(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n824_), .A2(new_n825_), .A3(new_n834_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n794_), .A2(new_n799_), .B1(new_n835_), .B2(new_n615_), .ZN(new_n836_));
  NOR4_X1   g635(.A1(new_n546_), .A2(new_n549_), .A3(new_n387_), .A4(new_n538_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G113gat), .B1(new_n839_), .B2(new_n626_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n830_), .A2(new_n319_), .A3(new_n833_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT57), .B1(new_n821_), .B2(new_n664_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT120), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n824_), .A2(new_n844_), .A3(new_n834_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n825_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n615_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n794_), .A2(new_n799_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n838_), .A2(KEYINPUT59), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT59), .B1(new_n836_), .B2(new_n838_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n626_), .A2(G113gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n840_), .B1(new_n853_), .B2(new_n854_), .ZN(G1340gat));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n746_), .A3(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G120gat), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT60), .ZN(new_n858_));
  AOI21_X1  g657(.A(G120gat), .B1(new_n746_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT121), .B1(new_n858_), .B2(G120gat), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n839_), .B(new_n861_), .C1(new_n859_), .C2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n857_), .A2(new_n863_), .ZN(G1341gat));
  AOI21_X1  g663(.A(G127gat), .B1(new_n839_), .B2(new_n616_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n616_), .A2(G127gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n853_), .B2(new_n866_), .ZN(G1342gat));
  INV_X1    g666(.A(new_n635_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G134gat), .B1(new_n839_), .B2(new_n868_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT122), .B(G134gat), .Z(new_n870_));
  NOR2_X1   g669(.A1(new_n318_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n853_), .B2(new_n871_), .ZN(G1343gat));
  NOR3_X1   g671(.A1(new_n527_), .A2(new_n549_), .A3(new_n548_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT123), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n836_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n626_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT124), .B(G141gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n746_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n835_), .A2(new_n615_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n848_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n874_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G155gat), .B1(new_n884_), .B2(new_n615_), .ZN(new_n885_));
  INV_X1    g684(.A(G155gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n876_), .A2(new_n886_), .A3(new_n616_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n885_), .A2(new_n889_), .A3(new_n887_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1346gat));
  AOI21_X1  g692(.A(G162gat), .B1(new_n876_), .B2(new_n868_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n675_), .A2(G162gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n876_), .B2(new_n895_), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n547_), .A2(new_n550_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n659_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n398_), .B1(new_n900_), .B2(new_n626_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n789_), .A2(new_n793_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n846_), .B2(new_n615_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n415_), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n903_), .A2(new_n904_), .A3(new_n625_), .A4(new_n899_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT62), .B1(new_n901_), .B2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n903_), .A2(new_n625_), .A3(new_n899_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n398_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n909_), .ZN(G1348gat));
  AOI21_X1  g709(.A(G176gat), .B1(new_n900_), .B2(new_n746_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n836_), .A2(new_n387_), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n897_), .A2(G176gat), .A3(new_n746_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1349gat));
  NAND3_X1  g713(.A1(new_n912_), .A2(new_n616_), .A3(new_n897_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n615_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n915_), .A2(new_n408_), .B1(new_n900_), .B2(new_n916_), .ZN(G1350gat));
  NAND2_X1  g716(.A1(new_n868_), .A2(new_n424_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT126), .Z(new_n919_));
  NAND2_X1  g718(.A1(new_n900_), .A2(new_n919_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n903_), .A2(new_n318_), .A3(new_n899_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n409_), .ZN(G1351gat));
  NOR3_X1   g721(.A1(new_n547_), .A2(new_n493_), .A3(new_n388_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n883_), .A2(new_n538_), .A3(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n625_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n351_), .ZN(G1352gat));
  OR2_X1    g725(.A1(new_n924_), .A2(new_n592_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(G204gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(new_n927_), .B2(new_n348_), .ZN(G1353gat));
  NOR2_X1   g728(.A1(new_n924_), .A2(new_n615_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n930_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT63), .B(G211gat), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n924_), .A2(new_n615_), .A3(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1354gat));
  INV_X1    g733(.A(new_n923_), .ZN(new_n935_));
  NOR4_X1   g734(.A1(new_n836_), .A2(new_n548_), .A3(new_n635_), .A4(new_n935_), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n319_), .A2(G218gat), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  OAI22_X1  g737(.A1(new_n936_), .A2(G218gat), .B1(new_n924_), .B2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  OAI221_X1 g740(.A(KEYINPUT127), .B1(new_n924_), .B2(new_n938_), .C1(new_n936_), .C2(G218gat), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1355gat));
endmodule


