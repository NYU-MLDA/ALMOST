//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT22), .B(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n207_), .B(KEYINPUT23), .Z(new_n208_));
  NOR2_X1   g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n206_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT26), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT26), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n213_), .A3(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n207_), .B(KEYINPUT23), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n202_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n216_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n210_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT85), .ZN(new_n224_));
  INV_X1    g023(.A(G197gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(G204gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT84), .B(G204gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(new_n225_), .ZN(new_n228_));
  INV_X1    g027(.A(G204gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT84), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT84), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G204gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n224_), .A3(G197gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT21), .B1(new_n228_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT21), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n225_), .A2(new_n229_), .ZN(new_n237_));
  AOI211_X1 g036(.A(new_n236_), .B(new_n237_), .C1(new_n233_), .C2(new_n225_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G211gat), .B(G218gat), .Z(new_n239_));
  NOR3_X1   g038(.A1(new_n235_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n228_), .A2(new_n234_), .A3(KEYINPUT21), .A4(new_n239_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n223_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT85), .B1(new_n229_), .B2(G197gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n244_), .B1(new_n233_), .B2(G197gat), .ZN(new_n245_));
  AOI211_X1 g044(.A(KEYINPUT85), .B(new_n225_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n236_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n237_), .B1(new_n233_), .B2(new_n225_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT21), .ZN(new_n249_));
  INV_X1    g048(.A(new_n239_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT78), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n214_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n212_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n213_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n221_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT79), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n219_), .A2(new_n220_), .ZN(new_n262_));
  OAI211_X1 g061(.A(KEYINPUT79), .B(new_n221_), .C1(new_n255_), .C2(new_n258_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(G183gat), .B1(new_n253_), .B2(new_n254_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n206_), .B1(new_n208_), .B2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n251_), .A2(new_n264_), .A3(new_n241_), .A4(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n243_), .A2(new_n267_), .A3(KEYINPUT20), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n251_), .A2(new_n241_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n264_), .A2(new_n266_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n210_), .A2(new_n222_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(new_n251_), .A3(new_n241_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n271_), .A3(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n273_), .A2(new_n280_), .A3(KEYINPUT87), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT87), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n277_), .A2(new_n282_), .A3(new_n271_), .A4(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G64gat), .B(G92gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n274_), .B1(new_n275_), .B2(new_n223_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(new_n271_), .A3(new_n267_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n271_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  AND4_X1   g094(.A1(KEYINPUT20), .A2(new_n243_), .A3(new_n267_), .A4(new_n271_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT91), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n289_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n290_), .B1(new_n298_), .B2(KEYINPUT92), .ZN(new_n299_));
  INV_X1    g098(.A(new_n289_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n264_), .A2(new_n266_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n228_), .A2(new_n234_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n239_), .B1(new_n302_), .B2(new_n236_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n242_), .B1(new_n303_), .B2(new_n249_), .ZN(new_n304_));
  OAI211_X1 g103(.A(KEYINPUT20), .B(new_n279_), .C1(new_n301_), .C2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n272_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n296_), .B1(new_n306_), .B2(KEYINPUT91), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n292_), .A2(new_n294_), .ZN(new_n308_));
  OAI211_X1 g107(.A(KEYINPUT92), .B(new_n300_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT27), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT93), .B1(new_n299_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n300_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n300_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT92), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT27), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(new_n298_), .B2(KEYINPUT92), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT93), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n281_), .A2(new_n283_), .A3(new_n300_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n320_), .A2(new_n312_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n311_), .A2(new_n319_), .B1(new_n316_), .B2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT81), .B(KEYINPUT2), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(G141gat), .B(G148gat), .C1(KEYINPUT81), .C2(KEYINPUT2), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n328_), .A2(KEYINPUT3), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n326_), .B(new_n327_), .C1(new_n329_), .C2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G155gat), .B(G162gat), .Z(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G155gat), .ZN(new_n336_));
  INV_X1    g135(.A(G162gat), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT1), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT1), .B1(new_n336_), .B2(new_n337_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n338_), .B(new_n339_), .C1(G155gat), .C2(G162gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(new_n325_), .A3(new_n330_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G127gat), .B(G134gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G113gat), .B(G120gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT89), .B1(new_n347_), .B2(KEYINPUT4), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n335_), .A2(new_n341_), .A3(new_n345_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(KEYINPUT4), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n342_), .A2(new_n353_), .A3(new_n354_), .A4(new_n346_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n348_), .A2(new_n350_), .A3(new_n352_), .A4(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n347_), .A2(new_n349_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n351_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G85gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT0), .B(G57gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n356_), .A2(new_n363_), .A3(new_n358_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n335_), .B2(new_n341_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n368_), .B1(new_n304_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n342_), .A2(KEYINPUT29), .ZN(new_n372_));
  INV_X1    g171(.A(new_n368_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n275_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(G228gat), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n371_), .A2(new_n374_), .A3(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(KEYINPUT82), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT28), .B1(new_n342_), .B2(KEYINPUT29), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT28), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n335_), .A2(new_n341_), .A3(new_n385_), .A4(new_n369_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G22gat), .B(G50gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n384_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n388_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n383_), .A2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n391_), .A2(new_n380_), .A3(KEYINPUT82), .A4(new_n382_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G15gat), .B(G43gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n345_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(new_n276_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(G71gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT30), .B(G99gat), .Z(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n398_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n395_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n405_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n367_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT90), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n366_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n366_), .A2(new_n411_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n363_), .B1(new_n357_), .B2(new_n352_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n348_), .A2(new_n355_), .A3(new_n350_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(new_n352_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n366_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n321_), .A2(new_n414_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n289_), .A2(KEYINPUT32), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n284_), .A2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n307_), .A2(new_n308_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n421_), .B(new_n367_), .C1(new_n422_), .C2(new_n420_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n395_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n323_), .A2(new_n409_), .B1(new_n424_), .B2(new_n405_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT75), .B(G15gat), .Z(new_n426_));
  INV_X1    g225(.A(G22gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G1gat), .ZN(new_n429_));
  INV_X1    g228(.A(G8gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT14), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT75), .B(G15gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(G22gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n428_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT76), .ZN(new_n435_));
  XOR2_X1   g234(.A(G1gat), .B(G8gat), .Z(new_n436_));
  INV_X1    g235(.A(KEYINPUT76), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n428_), .A2(new_n437_), .A3(new_n431_), .A4(new_n433_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n436_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G231gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT68), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G57gat), .B(G64gat), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(KEYINPUT11), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n446_), .A2(KEYINPUT11), .ZN(new_n449_));
  XOR2_X1   g248(.A(G71gat), .B(G78gat), .Z(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n445_), .A3(KEYINPUT11), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .A4(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(KEYINPUT11), .B2(new_n446_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n451_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(new_n447_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n456_), .B(KEYINPUT77), .Z(new_n457_));
  OR2_X1    g256(.A1(new_n444_), .A2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G127gat), .B(G155gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(G211gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT16), .B(G183gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n444_), .A2(new_n457_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n458_), .A2(KEYINPUT17), .A3(new_n462_), .A4(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n452_), .A2(KEYINPUT69), .A3(new_n455_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT69), .B1(new_n452_), .B2(new_n455_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n444_), .A2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n462_), .B(KEYINPUT17), .Z(new_n469_));
  NAND2_X1  g268(.A1(new_n444_), .A2(new_n467_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n464_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT74), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G85gat), .B(G92gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT66), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT7), .ZN(new_n478_));
  NOR2_X1   g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n475_), .B(KEYINPUT66), .C1(G99gat), .C2(G106gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n474_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT8), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT67), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT67), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n487_), .B1(new_n481_), .B2(new_n480_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n492_), .B(KEYINPUT8), .C1(new_n493_), .C2(new_n474_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT65), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n485_), .A2(new_n499_), .A3(new_n486_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  AOI211_X1 g300(.A(KEYINPUT8), .B(new_n474_), .C1(new_n501_), .C2(new_n482_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n495_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G29gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G85gat), .B(G92gat), .Z(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT9), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT9), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(G85gat), .A3(G92gat), .ZN(new_n511_));
  INV_X1    g310(.A(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(G99gat), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n513_), .A2(KEYINPUT10), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(KEYINPUT10), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n512_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n501_), .A2(new_n509_), .A3(new_n511_), .A4(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n504_), .A2(new_n507_), .A3(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n507_), .B(KEYINPUT15), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n502_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(KEYINPUT10), .B(G99gat), .Z(new_n523_));
  AOI22_X1  g322(.A1(new_n498_), .A2(new_n500_), .B1(new_n523_), .B2(new_n512_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n524_), .A2(KEYINPUT70), .A3(new_n509_), .A4(new_n511_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n519_), .B1(new_n520_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT34), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT35), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n529_), .A2(KEYINPUT35), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n518_), .A2(new_n527_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n530_), .B1(new_n518_), .B2(new_n527_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT73), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n518_), .A2(new_n527_), .A3(KEYINPUT73), .A4(new_n533_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n473_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(new_n337_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT72), .B(G134gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n518_), .A2(new_n527_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n536_), .B1(new_n545_), .B2(new_n531_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n534_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n538_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n544_), .B1(new_n548_), .B2(KEYINPUT36), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n543_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n539_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n539_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n551_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n550_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n553_), .B(new_n554_), .C1(new_n544_), .C2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n425_), .A2(new_n472_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n517_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n520_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n467_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G230gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT64), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n561_), .B2(new_n467_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n561_), .A2(new_n467_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT12), .B(new_n456_), .C1(new_n520_), .C2(new_n526_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n568_), .A2(new_n564_), .A3(new_n569_), .A4(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT5), .B(G176gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G204gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n566_), .A2(new_n571_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(KEYINPUT13), .A3(new_n579_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n507_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n441_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n507_), .A3(new_n439_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n585_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n519_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n589_), .A3(new_n585_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G169gat), .B(G197gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n591_), .A2(new_n593_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n593_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n599_), .B2(new_n590_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n584_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n559_), .A2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT94), .Z(new_n605_));
  INV_X1    g404(.A(new_n367_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608_));
  INV_X1    g407(.A(new_n538_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n519_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n522_), .A2(new_n525_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n504_), .B2(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n520_), .A2(new_n586_), .A3(new_n560_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n531_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT73), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n609_), .B1(new_n615_), .B2(new_n534_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n543_), .B1(new_n616_), .B2(new_n550_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n553_), .B1(new_n617_), .B2(new_n554_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n549_), .A2(new_n539_), .A3(new_n551_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n608_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n552_), .A2(new_n556_), .A3(KEYINPUT37), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n425_), .A2(new_n622_), .A3(new_n472_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(new_n603_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n429_), .A3(new_n367_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT38), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n607_), .A2(new_n626_), .ZN(G1324gat));
  INV_X1    g426(.A(new_n323_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n604_), .A2(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n629_), .A2(KEYINPUT96), .ZN(new_n630_));
  NAND2_X1  g429(.A1(KEYINPUT97), .A2(KEYINPUT39), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(KEYINPUT96), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n630_), .A2(G8gat), .A3(new_n631_), .A4(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(KEYINPUT97), .A2(KEYINPUT39), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n624_), .A2(new_n430_), .A3(new_n628_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT95), .Z(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n634_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n635_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(G1325gat));
  OAI21_X1  g440(.A(G15gat), .B1(new_n605_), .B2(new_n405_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT41), .Z(new_n643_));
  INV_X1    g442(.A(G15gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n624_), .A2(new_n644_), .A3(new_n407_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(G1326gat));
  INV_X1    g445(.A(new_n395_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G22gat), .B1(new_n605_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT42), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n624_), .A2(new_n427_), .A3(new_n395_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1327gat));
  INV_X1    g450(.A(new_n472_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n602_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(new_n425_), .A3(new_n557_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G29gat), .B1(new_n655_), .B2(new_n367_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n552_), .A2(new_n556_), .A3(KEYINPUT37), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT37), .B1(new_n552_), .B2(new_n556_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT43), .B1(new_n425_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n322_), .A2(new_n316_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n299_), .A2(new_n310_), .A3(KEYINPUT93), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n318_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n661_), .B(new_n409_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n419_), .A2(new_n423_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n405_), .A3(new_n647_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n622_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n654_), .B1(new_n660_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(KEYINPUT44), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n667_), .A2(new_n668_), .A3(new_n622_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n668_), .B1(new_n667_), .B2(new_n622_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n653_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT98), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n672_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(new_n606_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n670_), .A2(KEYINPUT44), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(G29gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n656_), .B1(new_n679_), .B2(new_n681_), .ZN(G1328gat));
  NOR2_X1   g481(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n323_), .B1(new_n670_), .B2(KEYINPUT44), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n684_), .B1(new_n672_), .B2(new_n677_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT99), .B(new_n684_), .C1(new_n672_), .C2(new_n677_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(G36gat), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n687_), .A2(KEYINPUT100), .A3(G36gat), .A4(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n655_), .A2(new_n694_), .A3(new_n628_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT45), .Z(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n683_), .B1(new_n693_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n683_), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n699_), .B(new_n696_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1329gat));
  NAND2_X1  g500(.A1(new_n680_), .A2(G43gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n678_), .A2(new_n702_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n703_), .A2(KEYINPUT102), .A3(new_n407_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT102), .B1(new_n703_), .B2(new_n407_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n655_), .A2(new_n407_), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n704_), .A2(new_n705_), .B1(G43gat), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n707_), .B(new_n709_), .ZN(G1330gat));
  AOI21_X1  g509(.A(G50gat), .B1(new_n655_), .B2(new_n395_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n678_), .A2(new_n647_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n680_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n584_), .A2(new_n601_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n623_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n367_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT104), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n559_), .A2(new_n715_), .ZN(new_n719_));
  INV_X1    g518(.A(G57gat), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n606_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1332gat));
  OAI21_X1  g521(.A(G64gat), .B1(new_n719_), .B2(new_n323_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n716_), .A2(new_n725_), .A3(new_n628_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n719_), .B2(new_n405_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  INV_X1    g528(.A(G71gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n716_), .A2(new_n730_), .A3(new_n407_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1334gat));
  OAI21_X1  g531(.A(G78gat), .B1(new_n719_), .B2(new_n647_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT105), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n716_), .A2(new_n395_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(G78gat), .B2(new_n736_), .ZN(G1335gat));
  NAND2_X1  g536(.A1(new_n715_), .A2(new_n472_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n738_), .A2(new_n425_), .A3(new_n557_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n367_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT106), .Z(new_n741_));
  AOI21_X1  g540(.A(new_n738_), .B1(new_n660_), .B2(new_n669_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n367_), .A2(G85gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n742_), .B2(new_n743_), .ZN(G1336gat));
  AOI21_X1  g543(.A(G92gat), .B1(new_n739_), .B2(new_n628_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n628_), .A2(G92gat), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT107), .Z(new_n747_));
  AOI21_X1  g546(.A(new_n745_), .B1(new_n742_), .B2(new_n747_), .ZN(G1337gat));
  AOI21_X1  g547(.A(new_n513_), .B1(new_n742_), .B2(new_n407_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n407_), .A2(new_n523_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n739_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(G1338gat));
  AOI21_X1  g552(.A(new_n512_), .B1(new_n742_), .B2(new_n395_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT52), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n739_), .A2(new_n512_), .A3(new_n395_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT109), .Z(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g558(.A(new_n585_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762_));
  OR3_X1    g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n597_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n592_), .A2(new_n589_), .A3(new_n760_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n761_), .B2(new_n597_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n580_), .A2(new_n598_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(new_n565_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n571_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n769_), .A2(new_n768_), .A3(new_n565_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n576_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT56), .B(new_n576_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n601_), .A2(new_n579_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT111), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n601_), .A2(new_n579_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n767_), .B1(new_n779_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(KEYINPUT57), .A4(new_n557_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n774_), .A2(new_n775_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n784_), .B1(new_n788_), .B2(new_n777_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n767_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT57), .B(new_n557_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT114), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n557_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n766_), .A2(new_n598_), .A3(new_n579_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT113), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n766_), .A2(new_n798_), .A3(new_n598_), .A4(new_n579_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n800_), .B(KEYINPUT58), .C1(new_n776_), .C2(new_n778_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n622_), .A3(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n787_), .A2(new_n792_), .A3(new_n795_), .A4(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n472_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n601_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n652_), .A2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT110), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n584_), .A3(new_n659_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT54), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n807_), .A2(new_n812_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n628_), .A2(new_n606_), .A3(new_n408_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816_), .B2(new_n601_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT115), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n806_), .A2(KEYINPUT116), .A3(new_n472_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT116), .B1(new_n806_), .B2(new_n472_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n812_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n823_), .A2(new_n814_), .B1(KEYINPUT59), .B2(new_n815_), .ZN(new_n824_));
  XOR2_X1   g623(.A(KEYINPUT117), .B(G113gat), .Z(new_n825_));
  NOR2_X1   g624(.A1(new_n808_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n818_), .B1(new_n824_), .B2(new_n826_), .ZN(G1340gat));
  INV_X1    g626(.A(G120gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n584_), .B2(KEYINPUT60), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n816_), .B(new_n829_), .C1(KEYINPUT60), .C2(new_n828_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n584_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n824_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n830_), .B1(new_n832_), .B2(new_n828_), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n816_), .B2(new_n652_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n824_), .A2(G127gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n652_), .ZN(G1342gat));
  AOI21_X1  g635(.A(G134gat), .B1(new_n816_), .B2(new_n558_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT118), .B(G134gat), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n659_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n824_), .B2(new_n839_), .ZN(G1343gat));
  AOI21_X1  g639(.A(new_n406_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n628_), .A2(new_n606_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n841_), .A2(KEYINPUT119), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT119), .B1(new_n841_), .B2(new_n842_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n601_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g645(.A(new_n831_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g647(.A(new_n652_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT120), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n851_), .B(new_n652_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT61), .B(G155gat), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n850_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1346gat));
  OAI21_X1  g655(.A(new_n622_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n337_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n558_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n337_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(KEYINPUT121), .A3(new_n337_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n858_), .B1(new_n862_), .B2(new_n863_), .ZN(G1347gat));
  NOR3_X1   g663(.A1(new_n323_), .A2(new_n367_), .A3(new_n408_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n821_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT124), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n821_), .A2(new_n868_), .A3(new_n865_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n601_), .A2(new_n204_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT125), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n323_), .A2(new_n367_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n601_), .A3(new_n407_), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT122), .Z(new_n876_));
  NAND3_X1  g675(.A1(new_n821_), .A2(new_n647_), .A3(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n821_), .A2(KEYINPUT123), .A3(new_n647_), .A4(new_n876_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(G169gat), .A3(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(KEYINPUT62), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(KEYINPUT62), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n873_), .B1(new_n882_), .B2(new_n883_), .ZN(G1348gat));
  AND4_X1   g683(.A1(G176gat), .A2(new_n813_), .A3(new_n831_), .A4(new_n865_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n870_), .A2(new_n831_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n205_), .ZN(G1349gat));
  NAND3_X1  g686(.A1(new_n813_), .A2(new_n652_), .A3(new_n865_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n888_), .A2(KEYINPUT126), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(KEYINPUT126), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n889_), .A2(new_n890_), .A3(G183gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n472_), .A2(new_n211_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n870_), .B2(new_n892_), .ZN(G1350gat));
  NAND4_X1  g692(.A1(new_n870_), .A2(new_n213_), .A3(new_n215_), .A4(new_n558_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n867_), .A2(new_n622_), .A3(new_n869_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n895_), .A2(new_n896_), .A3(G190gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n895_), .B2(G190gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n894_), .B1(new_n897_), .B2(new_n898_), .ZN(G1351gat));
  AND2_X1   g698(.A1(new_n841_), .A2(new_n874_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n601_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n831_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(G204gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(new_n227_), .B2(new_n903_), .ZN(G1353gat));
  NAND2_X1  g704(.A1(new_n900_), .A2(new_n652_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  AND2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n906_), .B2(new_n907_), .ZN(G1354gat));
  AOI21_X1  g709(.A(G218gat), .B1(new_n900_), .B2(new_n558_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n900_), .A2(new_n622_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(G218gat), .B2(new_n912_), .ZN(G1355gat));
endmodule


