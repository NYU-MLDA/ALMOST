//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_;
  AND2_X1   g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n203_));
  NOR2_X1   g002(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n205_), .B(new_n208_), .C1(G183gat), .C2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G169gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(G176gat), .B1(new_n211_), .B2(KEYINPUT76), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT22), .B(G169gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n212_), .B1(KEYINPUT76), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n209_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT75), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n206_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n202_), .A2(new_n207_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT74), .B(KEYINPUT23), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT75), .B1(new_n221_), .B2(new_n206_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT73), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT73), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(G169gat), .B2(G176gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT26), .B(G190gat), .ZN(new_n232_));
  INV_X1    g031(.A(G183gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT25), .B1(new_n233_), .B2(KEYINPUT72), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT72), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(G183gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n232_), .A2(new_n234_), .A3(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n226_), .A2(new_n228_), .A3(KEYINPUT24), .A4(new_n215_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n216_), .B1(new_n223_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G227gat), .A2(G233gat), .ZN(new_n242_));
  INV_X1    g041(.A(G15gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n241_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT77), .ZN(new_n247_));
  XOR2_X1   g046(.A(G127gat), .B(G134gat), .Z(new_n248_));
  INV_X1    g047(.A(G120gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G113gat), .ZN(new_n250_));
  INV_X1    g049(.A(G113gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G120gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n247_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n253_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G127gat), .B(G134gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n254_), .B1(new_n258_), .B2(new_n247_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n246_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G71gat), .B(G99gat), .ZN(new_n262_));
  INV_X1    g061(.A(G43gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT31), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n261_), .B(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G141gat), .ZN(new_n271_));
  INV_X1    g070(.A(G148gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT3), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT3), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(G141gat), .B2(G148gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT79), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n276_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n280_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n270_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT29), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT1), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(G155gat), .A3(G162gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n287_), .A3(new_n267_), .ZN(new_n288_));
  AND2_X1   g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT78), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n288_), .A2(KEYINPUT78), .A3(new_n291_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n283_), .A2(new_n284_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT28), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT28), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n283_), .A2(new_n296_), .A3(new_n299_), .A4(new_n284_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G22gat), .B(G50gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n298_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT81), .ZN(new_n306_));
  OAI22_X1  g105(.A1(new_n303_), .A2(new_n304_), .B1(KEYINPUT82), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n298_), .A2(new_n300_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n301_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n306_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n298_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n283_), .A2(new_n296_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT29), .ZN(new_n314_));
  OR2_X1    g113(.A1(G197gat), .A2(G204gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G197gat), .A2(G204gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(KEYINPUT21), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT21), .ZN(new_n318_));
  AND2_X1   g117(.A1(G197gat), .A2(G204gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G197gat), .A2(G204gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT80), .ZN(new_n324_));
  INV_X1    g123(.A(G218gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G211gat), .ZN(new_n326_));
  INV_X1    g125(.A(G211gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G218gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n329_), .A2(KEYINPUT21), .A3(new_n315_), .A4(new_n316_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n323_), .A2(new_n324_), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n324_), .B1(new_n323_), .B2(new_n330_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G228gat), .A2(G233gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n314_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n323_), .A2(new_n330_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n313_), .B2(KEYINPUT29), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n335_), .B1(new_n338_), .B2(new_n334_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n307_), .A2(new_n312_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n273_), .A2(new_n275_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT79), .B1(new_n342_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n276_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n269_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n288_), .A2(KEYINPUT78), .A3(new_n291_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT78), .B1(new_n288_), .B2(new_n291_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n259_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n283_), .A2(new_n258_), .A3(new_n296_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(KEYINPUT4), .A3(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT87), .B(KEYINPUT4), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n313_), .A2(new_n259_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G85gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT0), .B(G57gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n360_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n361_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n365_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n359_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n340_), .A2(new_n341_), .A3(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n374_));
  AND2_X1   g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT84), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT20), .B1(new_n333_), .B2(new_n241_), .ZN(new_n379_));
  OAI22_X1  g178(.A1(new_n220_), .A2(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n224_), .A2(KEYINPUT22), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n211_), .A2(new_n381_), .A3(new_n225_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT86), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n215_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n382_), .B2(new_n215_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n380_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT85), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n231_), .A2(new_n388_), .A3(new_n205_), .A4(new_n208_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n205_), .A2(new_n208_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT24), .B1(new_n226_), .B2(new_n228_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT85), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT25), .B(G183gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n232_), .A2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n394_), .A2(new_n239_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n389_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n337_), .B1(new_n387_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n378_), .B1(new_n379_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n333_), .A2(new_n241_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n387_), .A2(new_n396_), .A3(new_n337_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT20), .A4(new_n376_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G8gat), .B(G36gat), .Z(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT18), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n398_), .A2(new_n401_), .A3(new_n406_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT27), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(KEYINPUT92), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT92), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n398_), .A2(new_n414_), .A3(new_n401_), .A4(new_n406_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT93), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n387_), .A2(new_n396_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n336_), .ZN(new_n419_));
  OAI221_X1 g218(.A(new_n216_), .B1(new_n223_), .B2(new_n240_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(KEYINPUT20), .A4(new_n377_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT20), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(new_n376_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n411_), .B1(new_n423_), .B2(new_n407_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n416_), .A2(new_n417_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n417_), .B1(new_n416_), .B2(new_n424_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n373_), .B(new_n412_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n355_), .A2(new_n359_), .A3(new_n357_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n353_), .A2(new_n354_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n359_), .B1(new_n432_), .B2(KEYINPUT89), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n433_), .B1(KEYINPUT89), .B2(new_n432_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(new_n434_), .A3(new_n365_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT88), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n371_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT33), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n371_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n408_), .A2(new_n409_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n435_), .A2(new_n438_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n406_), .A2(KEYINPUT32), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n398_), .A2(new_n401_), .A3(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT91), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n423_), .A2(KEYINPUT32), .A3(new_n406_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n372_), .A3(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n340_), .A2(new_n341_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n427_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n340_), .A2(new_n341_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n412_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n266_), .A2(new_n372_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT94), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n412_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n416_), .A2(new_n424_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT93), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n416_), .A2(new_n417_), .A3(new_n424_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n456_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT94), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n451_), .A4(new_n453_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n266_), .A2(new_n450_), .B1(new_n455_), .B2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G85gat), .B(G92gat), .Z(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT10), .B(G99gat), .Z(new_n466_));
  INV_X1    g265(.A(G106gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G85gat), .ZN(new_n469_));
  INV_X1    g268(.A(G92gat), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT9), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G85gat), .B(G92gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT6), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n465_), .A2(new_n468_), .A3(new_n474_), .A4(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G57gat), .B(G64gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT11), .ZN(new_n479_));
  XOR2_X1   g278(.A(G71gat), .B(G78gat), .Z(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n478_), .A2(KEYINPUT11), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n480_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n475_), .B(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n464_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(KEYINPUT8), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n485_), .B(KEYINPUT7), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n472_), .B1(new_n492_), .B2(new_n476_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT8), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n477_), .B(new_n484_), .C1(new_n491_), .C2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT65), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n490_), .A2(KEYINPUT8), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n494_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n465_), .A2(new_n476_), .A3(new_n468_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n498_), .A2(new_n499_), .B1(new_n500_), .B2(new_n474_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT65), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n484_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n477_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n484_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n497_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(G230gat), .A2(G233gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n510_));
  NOR2_X1   g309(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n511_));
  OAI22_X1  g310(.A1(new_n501_), .A2(new_n484_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n508_), .B1(new_n501_), .B2(new_n484_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n511_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n504_), .A2(new_n505_), .A3(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G120gat), .B(G148gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT5), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G176gat), .B(G204gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n509_), .A2(new_n516_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT13), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n526_), .A2(KEYINPUT67), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(KEYINPUT67), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G1gat), .B(G8gat), .Z(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n533_));
  INV_X1    g332(.A(G1gat), .ZN(new_n534_));
  INV_X1    g333(.A(G8gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n533_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n531_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(new_n537_), .A3(new_n530_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G29gat), .B(G36gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n540_), .A2(new_n542_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n547_), .B(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n530_), .B1(new_n541_), .B2(new_n537_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n538_), .A2(new_n531_), .A3(new_n539_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n548_), .B(new_n549_), .C1(new_n551_), .C2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n549_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n548_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n547_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n555_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n463_), .A2(new_n529_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n501_), .A2(new_n547_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT34), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT35), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n570_), .B(new_n575_), .C1(new_n501_), .C2(new_n551_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n573_), .A2(new_n574_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n576_), .B(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G190gat), .B(G218gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n576_), .B(new_n577_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n584_), .B(KEYINPUT36), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT37), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n591_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n484_), .B(new_n596_), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(new_n554_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT17), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n598_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(KEYINPUT17), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n598_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n595_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n569_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n534_), .A3(new_n372_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT38), .ZN(new_n612_));
  INV_X1    g411(.A(new_n586_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n579_), .A2(new_n588_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n463_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n529_), .A2(new_n568_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n608_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT95), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(new_n372_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n612_), .B1(new_n534_), .B2(new_n621_), .ZN(G1324gat));
  INV_X1    g421(.A(new_n460_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n610_), .A2(new_n535_), .A3(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G8gat), .B1(new_n619_), .B2(new_n460_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n624_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI211_X1 g429(.A(KEYINPUT40), .B(new_n624_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1325gat));
  INV_X1    g431(.A(new_n266_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n610_), .A2(new_n243_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n620_), .A2(new_n633_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n635_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT41), .B1(new_n635_), .B2(G15gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(G1326gat));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n610_), .A2(new_n639_), .A3(new_n449_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT42), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n620_), .A2(new_n449_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(G22gat), .ZN(new_n643_));
  AOI211_X1 g442(.A(KEYINPUT42), .B(new_n639_), .C1(new_n620_), .C2(new_n449_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n643_), .B2(new_n644_), .ZN(G1327gat));
  NAND2_X1  g444(.A1(new_n615_), .A2(new_n608_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT96), .Z(new_n647_));
  NAND2_X1  g446(.A1(new_n569_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n372_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n594_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n592_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT43), .B1(new_n463_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n455_), .A2(new_n462_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n427_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n449_), .B1(new_n442_), .B2(new_n447_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n266_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(new_n595_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n653_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n527_), .A2(new_n528_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n608_), .A3(new_n567_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT44), .B1(new_n661_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  AOI211_X1 g465(.A(new_n666_), .B(new_n663_), .C1(new_n653_), .C2(new_n660_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n372_), .A2(G29gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n650_), .B1(new_n668_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(G36gat), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n569_), .A2(new_n671_), .A3(new_n623_), .A4(new_n647_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT45), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n665_), .A2(new_n667_), .A3(new_n460_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n671_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n673_), .B(KEYINPUT46), .C1(new_n674_), .C2(new_n671_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1329gat));
  AOI21_X1  g478(.A(new_n659_), .B1(new_n658_), .B2(new_n595_), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT43), .B(new_n652_), .C1(new_n654_), .C2(new_n657_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n664_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n666_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n664_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n266_), .A2(new_n263_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT97), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT97), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n683_), .A2(new_n684_), .A3(new_n688_), .A4(new_n685_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n263_), .B1(new_n648_), .B2(new_n266_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n687_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT47), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n687_), .A2(new_n693_), .A3(new_n689_), .A4(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1330gat));
  INV_X1    g494(.A(G50gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n649_), .A2(new_n696_), .A3(new_n449_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n668_), .A2(new_n449_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT98), .B1(new_n698_), .B2(G50gat), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT98), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n700_), .B(new_n696_), .C1(new_n668_), .C2(new_n449_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n699_), .B2(new_n701_), .ZN(G1331gat));
  NOR2_X1   g501(.A1(new_n608_), .A2(new_n567_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n616_), .A2(new_n529_), .A3(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT100), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(G57gat), .A3(new_n372_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT101), .ZN(new_n707_));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n529_), .A2(new_n609_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT99), .Z(new_n710_));
  NOR2_X1   g509(.A1(new_n463_), .A2(new_n567_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n372_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n708_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n707_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n706_), .A2(KEYINPUT101), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1332gat));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n705_), .A2(new_n623_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(G64gat), .ZN(new_n720_));
  INV_X1    g519(.A(G64gat), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT48), .B(new_n721_), .C1(new_n705_), .C2(new_n623_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n623_), .A2(new_n721_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT102), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n720_), .A2(new_n722_), .B1(new_n712_), .B2(new_n724_), .ZN(G1333gat));
  OR3_X1    g524(.A1(new_n712_), .A2(G71gat), .A3(new_n266_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n705_), .A2(new_n633_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT103), .B(KEYINPUT49), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(G71gat), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G71gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(G1334gat));
  INV_X1    g530(.A(KEYINPUT50), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n705_), .A2(new_n449_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G78gat), .ZN(new_n734_));
  INV_X1    g533(.A(G78gat), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT50), .B(new_n735_), .C1(new_n705_), .C2(new_n449_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n449_), .A2(new_n735_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT104), .Z(new_n738_));
  OAI22_X1  g537(.A1(new_n734_), .A2(new_n736_), .B1(new_n712_), .B2(new_n738_), .ZN(G1335gat));
  AND3_X1   g538(.A1(new_n711_), .A2(new_n529_), .A3(new_n647_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n469_), .A3(new_n372_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n527_), .A2(new_n608_), .A3(new_n568_), .A4(new_n528_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n661_), .A2(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(new_n372_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n741_), .B1(new_n746_), .B2(new_n469_), .ZN(G1336gat));
  NAND3_X1  g546(.A1(new_n745_), .A2(G92gat), .A3(new_n623_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n740_), .A2(new_n623_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n749_), .A2(KEYINPUT106), .A3(new_n470_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT106), .B1(new_n749_), .B2(new_n470_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT107), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n748_), .B(new_n754_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1337gat));
  NAND3_X1  g555(.A1(new_n740_), .A2(new_n466_), .A3(new_n633_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n745_), .A2(new_n633_), .ZN(new_n758_));
  INV_X1    g557(.A(G99gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n757_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT51), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(new_n757_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n740_), .A2(new_n467_), .A3(new_n449_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n661_), .A2(new_n744_), .A3(new_n449_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n765_), .B(new_n771_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1339gat));
  OAI21_X1  g574(.A(new_n703_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n525_), .B(KEYINPUT13), .Z(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT54), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n652_), .A2(new_n526_), .A3(new_n779_), .A4(new_n703_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n548_), .B(new_n556_), .C1(new_n551_), .C2(new_n554_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n549_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(new_n784_), .A3(new_n564_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n566_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n566_), .A2(new_n785_), .A3(KEYINPUT110), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n522_), .A2(new_n524_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n524_), .A2(new_n567_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n512_), .A2(new_n497_), .A3(new_n515_), .A4(new_n503_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n508_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n516_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT55), .A4(new_n515_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n521_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(KEYINPUT109), .A2(KEYINPUT56), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n791_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT109), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n797_), .A2(new_n802_), .A3(new_n803_), .A4(new_n521_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n790_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n782_), .B1(new_n805_), .B2(new_n615_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n512_), .A2(new_n515_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n808_), .A2(new_n513_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n788_), .A2(new_n789_), .B1(new_n809_), .B2(new_n523_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n797_), .A2(new_n803_), .A3(new_n521_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n803_), .B1(new_n797_), .B2(new_n521_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n807_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT58), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n807_), .B(new_n816_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n595_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n798_), .A2(new_n800_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n791_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n804_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n790_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n615_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n819_), .B1(new_n824_), .B2(KEYINPUT57), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n805_), .A2(KEYINPUT112), .A3(new_n782_), .A4(new_n615_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n806_), .B(new_n818_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n781_), .B1(new_n827_), .B2(new_n608_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n452_), .A2(new_n713_), .A3(new_n266_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n251_), .A3(new_n567_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n818_), .A2(new_n806_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT113), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n824_), .A2(KEYINPUT57), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT112), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n824_), .A2(new_n819_), .A3(KEYINPUT57), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n818_), .A2(new_n839_), .A3(new_n806_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n834_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n781_), .B1(new_n841_), .B2(new_n608_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n830_), .A2(KEYINPUT59), .ZN(new_n844_));
  INV_X1    g643(.A(new_n831_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n843_), .A2(new_n844_), .B1(new_n845_), .B2(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n567_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n832_), .B1(new_n848_), .B2(new_n251_), .ZN(G1340gat));
  OAI21_X1  g648(.A(KEYINPUT59), .B1(new_n828_), .B2(new_n830_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n844_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n850_), .B(new_n529_), .C1(new_n842_), .C2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n249_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n853_), .B2(new_n852_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n249_), .B1(new_n662_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n831_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n249_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1341gat));
  AOI21_X1  g657(.A(G127gat), .B1(new_n831_), .B2(new_n618_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n618_), .A2(G127gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT115), .Z(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n846_), .B2(new_n861_), .ZN(G1342gat));
  OAI211_X1 g661(.A(new_n850_), .B(new_n595_), .C1(new_n842_), .C2(new_n851_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G134gat), .ZN(new_n864_));
  INV_X1    g663(.A(G134gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n831_), .A2(new_n865_), .A3(new_n615_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n864_), .A2(KEYINPUT116), .A3(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1343gat));
  NAND2_X1  g670(.A1(new_n827_), .A2(new_n608_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n781_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n460_), .A2(new_n372_), .A3(new_n266_), .A4(new_n449_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT117), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n874_), .A2(KEYINPUT118), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(KEYINPUT118), .B1(new_n874_), .B2(new_n876_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n567_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g679(.A(new_n529_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g681(.A(new_n618_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  NOR2_X1   g684(.A1(new_n877_), .A2(new_n878_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G162gat), .B1(new_n886_), .B2(new_n652_), .ZN(new_n887_));
  INV_X1    g686(.A(G162gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n615_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n886_), .B2(new_n889_), .ZN(G1347gat));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n623_), .A2(new_n453_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n449_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n833_), .A2(KEYINPUT113), .B1(new_n836_), .B2(new_n837_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n618_), .B1(new_n894_), .B2(new_n840_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n567_), .B(new_n893_), .C1(new_n895_), .C2(new_n781_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n843_), .A2(new_n213_), .A3(new_n567_), .A4(new_n893_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT62), .B1(new_n896_), .B2(G169gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n891_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n896_), .A2(G169gat), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n904_), .A2(KEYINPUT119), .A3(new_n898_), .A4(new_n897_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n901_), .A2(new_n905_), .ZN(G1348gat));
  NAND2_X1  g705(.A1(new_n843_), .A2(new_n893_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G176gat), .B1(new_n908_), .B2(new_n529_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n828_), .A2(new_n449_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n662_), .A2(new_n225_), .A3(new_n892_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(G1349gat));
  NAND4_X1  g711(.A1(new_n910_), .A2(new_n623_), .A3(new_n453_), .A4(new_n618_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n233_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n608_), .A2(new_n393_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n907_), .B2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(KEYINPUT120), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n914_), .B(new_n918_), .C1(new_n907_), .C2(new_n915_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n907_), .B2(new_n652_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n615_), .A2(new_n232_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n907_), .B2(new_n922_), .ZN(G1351gat));
  AND2_X1   g722(.A1(new_n373_), .A2(new_n266_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n623_), .A2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(KEYINPUT121), .B1(new_n874_), .B2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n828_), .A2(new_n928_), .A3(new_n925_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(G197gat), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n930_), .A2(new_n568_), .A3(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n930_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n567_), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT122), .B(G197gat), .Z(new_n936_));
  AOI21_X1  g735(.A(new_n933_), .B1(new_n935_), .B2(new_n936_), .ZN(G1352gat));
  NOR2_X1   g736(.A1(new_n930_), .A2(new_n662_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(KEYINPUT123), .B(G204gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n938_), .B(new_n939_), .ZN(G1353gat));
  AOI21_X1  g739(.A(new_n608_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n934_), .A2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(KEYINPUT124), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n942_), .A2(new_n945_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n934_), .A2(new_n944_), .A3(new_n941_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1354gat));
  XOR2_X1   g747(.A(KEYINPUT126), .B(G218gat), .Z(new_n949_));
  NOR2_X1   g748(.A1(new_n652_), .A2(new_n949_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(KEYINPUT127), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n930_), .A2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n953_));
  INV_X1    g752(.A(new_n615_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n930_), .B2(new_n954_), .ZN(new_n955_));
  OAI211_X1 g754(.A(KEYINPUT125), .B(new_n615_), .C1(new_n927_), .C2(new_n929_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n955_), .A2(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n952_), .B1(new_n957_), .B2(new_n949_), .ZN(G1355gat));
endmodule


