//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n909_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT36), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT10), .B(G99gat), .Z(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT9), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n216_));
  INV_X1    g015(.A(G85gat), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n214_), .A2(new_n215_), .A3(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n215_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n208_), .B(new_n211_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n224_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT7), .ZN(new_n229_));
  INV_X1    g028(.A(G99gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n210_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(KEYINPUT66), .A3(new_n225_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n208_), .A3(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n212_), .A2(new_n213_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n223_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT65), .B(KEYINPUT8), .Z(new_n237_));
  NOR2_X1   g036(.A1(new_n226_), .A2(new_n227_), .ZN(new_n238_));
  AOI211_X1 g037(.A(new_n237_), .B(new_n234_), .C1(new_n208_), .C2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n222_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G29gat), .B(G36gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G43gat), .B(G50gat), .Z(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n241_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT15), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n240_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n240_), .A2(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n222_), .B(KEYINPUT67), .C1(new_n236_), .C2(new_n239_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n247_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n251_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(KEYINPUT73), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G232gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT34), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(KEYINPUT35), .A3(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(KEYINPUT35), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT72), .Z(new_n263_));
  AND3_X1   g062(.A1(new_n257_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n261_), .B1(new_n257_), .B2(new_n263_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n206_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT74), .B1(new_n264_), .B2(new_n265_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n204_), .A2(new_n205_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n268_), .ZN(new_n270_));
  OAI221_X1 g069(.A(KEYINPUT74), .B1(new_n270_), .B2(new_n206_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G127gat), .B(G155gat), .ZN(new_n279_));
  INV_X1    g078(.A(G211gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(KEYINPUT16), .B(G183gat), .Z(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G57gat), .B(G64gat), .Z(new_n285_));
  INV_X1    g084(.A(KEYINPUT11), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G71gat), .B(G78gat), .Z(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT68), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n285_), .A2(new_n286_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n287_), .A2(new_n292_), .A3(new_n288_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n290_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n291_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G231gat), .ZN(new_n297_));
  INV_X1    g096(.A(G233gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n296_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G15gat), .B(G22gat), .ZN(new_n301_));
  INV_X1    g100(.A(G1gat), .ZN(new_n302_));
  INV_X1    g101(.A(G8gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT14), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G1gat), .B(G8gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n300_), .B(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n284_), .B1(new_n309_), .B2(KEYINPUT76), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT17), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n284_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT17), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n278_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT77), .ZN(new_n318_));
  OR2_X1    g117(.A1(G113gat), .A2(G120gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G113gat), .A2(G120gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G127gat), .ZN(new_n322_));
  INV_X1    g121(.A(G134gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G127gat), .A2(G134gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT83), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT83), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n321_), .A2(new_n326_), .A3(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n319_), .A2(new_n324_), .A3(new_n325_), .A4(new_n320_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n331_), .A2(KEYINPUT84), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(KEYINPUT84), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n328_), .B(new_n330_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G155gat), .ZN(new_n336_));
  INV_X1    g135(.A(G162gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT1), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G155gat), .A3(G162gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(new_n337_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(G141gat), .ZN(new_n344_));
  INV_X1    g143(.A(G148gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT2), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n343_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n349_), .A2(new_n351_), .A3(new_n352_), .A4(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G155gat), .B(G162gat), .Z(new_n355_));
  AND3_X1   g154(.A1(new_n354_), .A2(KEYINPUT86), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT86), .B1(new_n354_), .B2(new_n355_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n347_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n335_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n327_), .A2(new_n331_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n347_), .B(new_n361_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n342_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n354_), .A2(new_n355_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n354_), .A2(KEYINPUT86), .A3(new_n355_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n365_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(KEYINPUT4), .B(new_n362_), .C1(new_n370_), .C2(new_n334_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n335_), .A2(new_n372_), .A3(new_n358_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n373_), .A3(KEYINPUT100), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT100), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n359_), .A2(new_n375_), .A3(KEYINPUT4), .A4(new_n362_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n360_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n364_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT101), .B(KEYINPUT0), .Z(new_n380_));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT33), .B1(new_n379_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n360_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388_));
  NOR4_X1   g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n384_), .A4(new_n364_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n378_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n359_), .A2(new_n378_), .A3(new_n362_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n384_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT99), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G197gat), .B(G204gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT21), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT91), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT92), .ZN(new_n403_));
  INV_X1    g202(.A(G197gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(G204gat), .ZN(new_n405_));
  INV_X1    g204(.A(G204gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT92), .B1(new_n406_), .B2(G197gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(G197gat), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n401_), .B(new_n405_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n404_), .A2(G204gat), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n410_), .B(KEYINPUT21), .C1(new_n408_), .C2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G218gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n280_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G211gat), .A2(G218gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n402_), .A2(new_n409_), .A3(new_n412_), .A4(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT93), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n405_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n414_), .A2(KEYINPUT93), .A3(new_n415_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(KEYINPUT21), .A4(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT26), .B(G190gat), .ZN(new_n425_));
  INV_X1    g224(.A(G183gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT25), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT25), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n426_), .B2(KEYINPUT25), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n425_), .A2(new_n427_), .A3(new_n429_), .A4(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT24), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n433_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G183gat), .A2(G190gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT23), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444_));
  INV_X1    g243(.A(G169gat), .ZN(new_n445_));
  INV_X1    g244(.A(G176gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G169gat), .A2(G176gat), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n447_), .A2(KEYINPUT24), .A3(new_n448_), .A4(new_n434_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n432_), .A2(new_n437_), .A3(new_n443_), .A4(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(G183gat), .A2(G190gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n440_), .A2(new_n451_), .A3(new_n441_), .ZN(new_n452_));
  AND2_X1   g251(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n446_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n455_), .A3(new_n448_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n399_), .B1(new_n424_), .B2(new_n457_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n453_), .A2(new_n454_), .A3(KEYINPUT96), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT96), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT22), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n445_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n460_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n446_), .B1(new_n459_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n452_), .A2(new_n448_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT97), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT96), .B1(new_n453_), .B2(new_n454_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n462_), .A2(new_n460_), .A3(new_n463_), .ZN(new_n470_));
  AOI21_X1  g269(.A(G176gat), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n452_), .A2(new_n448_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT97), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT25), .B(G183gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n442_), .B1(new_n474_), .B2(new_n425_), .ZN(new_n475_));
  AND2_X1   g274(.A1(KEYINPUT95), .A2(KEYINPUT24), .ZN(new_n476_));
  NOR2_X1   g275(.A1(KEYINPUT95), .A2(KEYINPUT24), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n478_), .A2(new_n448_), .A3(new_n447_), .A4(new_n434_), .ZN(new_n479_));
  OAI22_X1  g278(.A1(new_n435_), .A2(new_n436_), .B1(new_n477_), .B2(new_n476_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n475_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n468_), .A2(new_n473_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n423_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n398_), .B1(new_n458_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n450_), .A2(new_n456_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n423_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(KEYINPUT20), .A3(new_n398_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n482_), .A2(new_n423_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT98), .B(KEYINPUT18), .Z(new_n490_));
  XNOR2_X1  g289(.A(G8gat), .B(G36gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G64gat), .B(G92gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n484_), .A2(new_n489_), .A3(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n482_), .A2(new_n423_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT20), .B1(new_n423_), .B2(new_n485_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n397_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n399_), .B1(new_n423_), .B2(new_n485_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n500_), .B(new_n398_), .C1(new_n423_), .C2(new_n482_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n494_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n395_), .B1(new_n496_), .B2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n495_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n494_), .A3(new_n501_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT99), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n394_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n377_), .A2(new_n378_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(new_n385_), .A3(new_n363_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n384_), .B1(new_n387_), .B2(new_n364_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n458_), .A2(new_n398_), .A3(new_n483_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n465_), .A2(new_n466_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n481_), .A2(new_n512_), .A3(new_n422_), .A4(new_n417_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n486_), .A2(new_n513_), .A3(KEYINPUT20), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n397_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n494_), .A2(KEYINPUT32), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n509_), .A2(new_n510_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n484_), .A2(new_n489_), .A3(new_n517_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n390_), .A2(new_n507_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G22gat), .B(G50gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT87), .ZN(new_n522_));
  XOR2_X1   g321(.A(G78gat), .B(G106gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n526_), .A2(G228gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(G228gat), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n298_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n529_), .B(KEYINPUT90), .Z(new_n530_));
  NAND3_X1  g329(.A1(new_n358_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n423_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT88), .B1(new_n358_), .B2(KEYINPUT29), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n530_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n530_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n358_), .A2(KEYINPUT94), .A3(KEYINPUT29), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT94), .B1(new_n358_), .B2(KEYINPUT29), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n535_), .B(new_n423_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  OR3_X1    g337(.A1(new_n358_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT28), .B1(new_n358_), .B2(KEYINPUT29), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n534_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n534_), .B2(new_n538_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n525_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n534_), .A2(new_n538_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n541_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n534_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n524_), .A3(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n544_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n544_), .A2(new_n549_), .A3(new_n510_), .A4(new_n509_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n516_), .A2(new_n495_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(KEYINPUT27), .A3(new_n505_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT102), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT27), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n496_), .B2(new_n502_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n516_), .B2(new_n495_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT102), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n505_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n554_), .A2(new_n556_), .A3(new_n559_), .ZN(new_n560_));
  OAI22_X1  g359(.A1(new_n520_), .A2(new_n550_), .B1(new_n551_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G15gat), .B(G43gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(new_n230_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT30), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n457_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT82), .B(G71gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G227gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n565_), .A2(new_n569_), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n570_), .A2(new_n571_), .A3(KEYINPUT85), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n334_), .B(KEYINPUT31), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n572_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT103), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n560_), .B2(new_n550_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n557_), .A2(new_n558_), .A3(new_n505_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n558_), .B1(new_n557_), .B2(new_n505_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n544_), .A2(new_n549_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n580_), .A2(KEYINPUT103), .A3(new_n581_), .A4(new_n556_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n509_), .A2(new_n510_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n575_), .A2(new_n584_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n561_), .A2(new_n575_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT78), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n307_), .A2(new_n247_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n249_), .B2(new_n307_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n307_), .B(new_n247_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n590_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n587_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n587_), .B2(new_n594_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT79), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G169gat), .B(G197gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n598_), .B(new_n599_), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n596_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT71), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n294_), .A2(new_n295_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n255_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n296_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n606_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n296_), .A2(KEYINPUT12), .A3(new_n240_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n613_), .A2(new_n605_), .A3(new_n608_), .A4(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(KEYINPUT5), .B(G176gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT70), .B(G204gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n610_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n603_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n610_), .A2(new_n615_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n620_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n610_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(KEYINPUT71), .A3(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n624_), .A2(new_n628_), .A3(KEYINPUT13), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT13), .B1(new_n624_), .B2(new_n628_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n586_), .A2(new_n602_), .A3(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n318_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n302_), .A3(new_n584_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT38), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n315_), .A2(new_n272_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n584_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G1gat), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(G1324gat));
  NAND3_X1  g439(.A1(new_n633_), .A2(new_n303_), .A3(new_n560_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n560_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G8gat), .B1(new_n637_), .B2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(KEYINPUT39), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(KEYINPUT39), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n646_), .B(new_n647_), .Z(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n637_), .B2(new_n575_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT105), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n575_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n633_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n652_), .B(new_n653_), .C1(G15gat), .C2(new_n655_), .ZN(G1326gat));
  OAI21_X1  g455(.A(G22gat), .B1(new_n637_), .B2(new_n581_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT42), .ZN(new_n658_));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n633_), .A2(new_n659_), .A3(new_n550_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(G1327gat));
  NOR2_X1   g460(.A1(new_n631_), .A2(new_n602_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n663_));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n269_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n273_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n275_), .A2(KEYINPUT107), .A3(new_n276_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n583_), .A2(new_n585_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n503_), .A2(new_n506_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n394_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n509_), .A2(new_n388_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n379_), .A2(KEYINPUT33), .A3(new_n385_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n671_), .A2(new_n672_), .A3(new_n673_), .A4(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n518_), .A2(new_n519_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n550_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n560_), .A2(new_n551_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n575_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n670_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n663_), .B1(new_n669_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n277_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n586_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n315_), .B(new_n662_), .C1(new_n681_), .C2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT43), .B1(new_n275_), .B2(new_n276_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n680_), .A2(new_n688_), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n668_), .A2(new_n667_), .B1(new_n670_), .B2(new_n679_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(new_n663_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n691_), .A2(KEYINPUT44), .A3(new_n315_), .A4(new_n662_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n687_), .A2(G29gat), .A3(new_n584_), .A4(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n315_), .A2(new_n272_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n632_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(new_n638_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(G29gat), .B2(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT108), .Z(G1328gat));
  OR2_X1    g498(.A1(new_n642_), .A2(KEYINPUT109), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n642_), .A2(KEYINPUT109), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n696_), .A2(G36gat), .A3(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT45), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n687_), .A2(new_n560_), .A3(new_n692_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n704_), .A2(KEYINPUT46), .A3(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1329gat));
  INV_X1    g510(.A(G43gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(new_n696_), .B2(new_n575_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n575_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n714_));
  AND4_X1   g513(.A1(KEYINPUT110), .A2(new_n714_), .A3(G43gat), .A4(new_n692_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n692_), .A2(G43gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT110), .B1(new_n716_), .B2(new_n714_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n713_), .B(new_n719_), .C1(new_n715_), .C2(new_n717_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1330gat));
  INV_X1    g522(.A(new_n696_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G50gat), .B1(new_n724_), .B2(new_n550_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n687_), .A2(G50gat), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n692_), .A2(new_n550_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n726_), .B2(new_n727_), .ZN(G1331gat));
  NAND2_X1  g527(.A1(new_n624_), .A2(new_n628_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT13), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n624_), .A2(new_n628_), .A3(KEYINPUT13), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n602_), .A3(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n586_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n636_), .ZN(new_n735_));
  INV_X1    g534(.A(G57gat), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n638_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n318_), .A2(new_n734_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n638_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(new_n739_), .B2(new_n738_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n737_), .B1(new_n741_), .B2(new_n736_), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n735_), .B2(new_n702_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(G64gat), .ZN(new_n746_));
  INV_X1    g545(.A(new_n702_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n738_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1333gat));
  OAI21_X1  g548(.A(G71gat), .B1(new_n735_), .B2(new_n575_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT49), .ZN(new_n751_));
  INV_X1    g550(.A(G71gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n738_), .A2(new_n752_), .A3(new_n654_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1334gat));
  OAI21_X1  g553(.A(G78gat), .B1(new_n735_), .B2(new_n581_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT50), .ZN(new_n756_));
  INV_X1    g555(.A(G78gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n738_), .A2(new_n757_), .A3(new_n550_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1335gat));
  NOR3_X1   g558(.A1(new_n586_), .A2(new_n694_), .A3(new_n733_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n761_), .A2(G85gat), .A3(new_n638_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n733_), .B2(new_n316_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n631_), .A2(KEYINPUT114), .A3(new_n315_), .A4(new_n602_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n691_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n584_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n762_), .B1(new_n768_), .B2(G85gat), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT115), .Z(G1336gat));
  NAND3_X1  g569(.A1(new_n767_), .A2(G92gat), .A3(new_n747_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n218_), .B1(new_n761_), .B2(new_n642_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT116), .ZN(G1337gat));
  NAND4_X1  g573(.A1(new_n760_), .A2(KEYINPUT117), .A3(new_n209_), .A4(new_n654_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n629_), .A2(new_n630_), .A3(new_n601_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n680_), .A2(new_n209_), .A3(new_n695_), .A4(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n778_), .B2(new_n575_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n775_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n766_), .B(new_n654_), .C1(new_n681_), .C2(new_n684_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G99gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n782_), .A3(KEYINPUT119), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n780_), .A2(new_n782_), .A3(KEYINPUT118), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT51), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n789_), .A2(KEYINPUT51), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n783_), .A2(new_n784_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT120), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n794_), .B2(new_n786_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n791_), .A2(new_n795_), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n760_), .A2(new_n210_), .A3(new_n550_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n767_), .A2(new_n550_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(G106gat), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT52), .B(new_n210_), .C1(new_n767_), .C2(new_n550_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g602(.A1(new_n316_), .A2(new_n275_), .A3(new_n602_), .A4(new_n276_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n631_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(KEYINPUT121), .A2(KEYINPUT54), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n805_), .A2(new_n806_), .A3(new_n809_), .A4(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n807_), .B(new_n808_), .C1(new_n804_), .C2(new_n631_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n613_), .A2(new_n605_), .A3(new_n614_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n609_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n615_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n815_), .A2(new_n814_), .A3(new_n609_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n620_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT56), .B(new_n620_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n592_), .A2(new_n590_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n600_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n596_), .A2(new_n600_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(new_n627_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n824_), .A2(KEYINPUT58), .A3(new_n627_), .A4(new_n827_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n277_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n272_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n601_), .A2(new_n627_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n624_), .A2(new_n628_), .A3(new_n827_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n833_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT57), .B(new_n833_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n832_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n813_), .B1(new_n841_), .B2(new_n315_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n583_), .A2(new_n584_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n842_), .A2(new_n575_), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n601_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n841_), .A2(new_n315_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n813_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n575_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n843_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n846_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n842_), .A2(KEYINPUT59), .A3(new_n575_), .A4(new_n843_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n602_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n845_), .B1(new_n853_), .B2(G113gat), .ZN(G1340gat));
  NOR3_X1   g653(.A1(new_n851_), .A2(new_n852_), .A3(new_n806_), .ZN(new_n855_));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(KEYINPUT60), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n842_), .A2(new_n575_), .A3(new_n843_), .A4(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n806_), .B2(KEYINPUT60), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n855_), .A2(new_n856_), .B1(new_n861_), .B2(new_n862_), .ZN(G1341gat));
  AOI21_X1  g662(.A(G127gat), .B1(new_n844_), .B2(new_n316_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n851_), .A2(new_n852_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n315_), .A2(new_n322_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(G1342gat));
  AOI21_X1  g666(.A(G134gat), .B1(new_n844_), .B2(new_n272_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n278_), .A2(new_n323_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n865_), .B2(new_n869_), .ZN(G1343gat));
  NOR2_X1   g669(.A1(new_n842_), .A2(new_n654_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n747_), .A2(new_n638_), .A3(new_n581_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n344_), .A3(new_n601_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G141gat), .B1(new_n873_), .B2(new_n602_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1344gat));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n345_), .A3(new_n631_), .ZN(new_n878_));
  OAI21_X1  g677(.A(G148gat), .B1(new_n873_), .B2(new_n806_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1345gat));
  NAND3_X1  g679(.A1(new_n871_), .A2(new_n316_), .A3(new_n872_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  INV_X1    g682(.A(new_n669_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n873_), .A2(new_n337_), .A3(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n847_), .A2(new_n848_), .ZN(new_n887_));
  AND4_X1   g686(.A1(new_n272_), .A2(new_n887_), .A3(new_n575_), .A4(new_n872_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n886_), .B1(new_n888_), .B2(G162gat), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT123), .B(new_n337_), .C1(new_n873_), .C2(new_n833_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n885_), .B1(new_n889_), .B2(new_n890_), .ZN(G1347gat));
  XNOR2_X1  g690(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n842_), .A2(new_n584_), .A3(new_n575_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n702_), .A2(new_n550_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  OAI211_X1 g694(.A(G169gat), .B(new_n892_), .C1(new_n895_), .C2(new_n602_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n892_), .ZN(new_n897_));
  AND4_X1   g696(.A1(new_n601_), .A2(new_n887_), .A3(new_n585_), .A4(new_n894_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n445_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n464_), .B2(new_n459_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n896_), .A2(new_n899_), .A3(new_n900_), .ZN(G1348gat));
  NAND3_X1  g700(.A1(new_n893_), .A2(new_n631_), .A3(new_n894_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g702(.A1(new_n887_), .A2(new_n316_), .A3(new_n585_), .A4(new_n894_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n474_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n426_), .B2(new_n904_), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n895_), .B2(new_n278_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n272_), .A2(new_n425_), .ZN(new_n908_));
  XOR2_X1   g707(.A(new_n908_), .B(KEYINPUT125), .Z(new_n909_));
  OAI21_X1  g708(.A(new_n907_), .B1(new_n895_), .B2(new_n909_), .ZN(G1351gat));
  NOR3_X1   g709(.A1(new_n842_), .A2(new_n551_), .A3(new_n654_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n601_), .A3(new_n747_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g712(.A1(new_n911_), .A2(new_n631_), .A3(new_n747_), .ZN(new_n914_));
  AND2_X1   g713(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n915_));
  NOR2_X1   g714(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n914_), .B2(new_n915_), .ZN(G1353gat));
  AOI21_X1  g717(.A(new_n315_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT127), .Z(new_n920_));
  NAND3_X1  g719(.A1(new_n911_), .A2(new_n747_), .A3(new_n920_), .ZN(new_n921_));
  OR2_X1    g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1354gat));
  AND4_X1   g722(.A1(G218gat), .A2(new_n911_), .A3(new_n277_), .A4(new_n747_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n911_), .A2(new_n272_), .A3(new_n747_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n413_), .B2(new_n925_), .ZN(G1355gat));
endmodule


