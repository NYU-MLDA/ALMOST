//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n202_), .A2(new_n203_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(KEYINPUT15), .A3(new_n205_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT77), .B(G8gat), .Z(new_n211_));
  INV_X1    g010(.A(G1gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT76), .B(G15gat), .ZN(new_n214_));
  INV_X1    g013(.A(G22gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n215_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G1gat), .B(G8gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n220_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n210_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT81), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT81), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n210_), .A2(new_n221_), .A3(new_n225_), .A4(new_n222_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n221_), .A2(new_n222_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n230_), .B2(new_n206_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n206_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n221_), .A2(new_n205_), .A3(new_n204_), .A4(new_n222_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n229_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G169gat), .B(G197gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  AND3_X1   g038(.A1(new_n232_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G226gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT19), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(G183gat), .A3(G190gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G183gat), .ZN(new_n249_));
  INV_X1    g048(.A(G190gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT23), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n248_), .B(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT82), .B(G176gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT22), .B(G169gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(KEYINPUT83), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n258_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT83), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n255_), .A2(new_n256_), .A3(new_n259_), .A4(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT24), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n264_), .A2(KEYINPUT24), .A3(new_n256_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT25), .B(G183gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G190gat), .ZN(new_n268_));
  AOI211_X1 g067(.A(new_n265_), .B(new_n266_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n251_), .A2(new_n246_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G211gat), .B(G218gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT91), .Z(new_n274_));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT21), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n273_), .B(KEYINPUT91), .ZN(new_n279_));
  INV_X1    g078(.A(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n276_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT20), .B1(new_n272_), .B2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n278_), .A2(new_n282_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n260_), .A2(new_n256_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT96), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n286_), .A2(new_n287_), .B1(new_n270_), .B2(new_n254_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(new_n287_), .B2(new_n286_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n269_), .A2(new_n252_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OAI22_X1  g090(.A1(new_n284_), .A2(KEYINPUT95), .B1(new_n285_), .B2(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n284_), .A2(KEYINPUT95), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n244_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n285_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n272_), .A2(new_n283_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n295_), .A2(KEYINPUT20), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n244_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G8gat), .B(G36gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT18), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G64gat), .B(G92gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n294_), .A2(new_n304_), .A3(new_n299_), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT27), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(KEYINPUT100), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n297_), .A2(new_n298_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n292_), .A2(new_n293_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(new_n298_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n312_), .A2(new_n304_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(KEYINPUT100), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n309_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n308_), .B1(new_n315_), .B2(KEYINPUT27), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G225gat), .A2(G233gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G141gat), .A2(G148gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(G155gat), .A3(G162gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT89), .Z(new_n324_));
  INV_X1    g123(.A(G155gat), .ZN(new_n325_));
  INV_X1    g124(.A(G162gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(KEYINPUT88), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT88), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(G155gat), .B2(G162gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n322_), .B1(G155gat), .B2(G162gat), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n319_), .B(new_n321_), .C1(new_n324_), .C2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n330_), .B1(G155gat), .B2(G162gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n320_), .B(KEYINPUT3), .Z(new_n335_));
  XOR2_X1   g134(.A(new_n319_), .B(KEYINPUT2), .Z(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G127gat), .B(G134gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n333_), .A2(new_n337_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n318_), .B1(new_n342_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT4), .B1(new_n343_), .B2(new_n346_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n342_), .A2(new_n347_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(KEYINPUT4), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n348_), .B1(new_n351_), .B2(new_n318_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G57gat), .B(G85gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n352_), .B(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n358_), .B(KEYINPUT99), .Z(new_n359_));
  XNOR2_X1  g158(.A(new_n346_), .B(KEYINPUT31), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362_));
  INV_X1    g161(.A(G43gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365_));
  INV_X1    g164(.A(G15gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n364_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n272_), .B(KEYINPUT30), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT85), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n370_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n368_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n368_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n361_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n368_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n372_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n369_), .A2(new_n370_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(new_n374_), .A3(new_n360_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n376_), .A2(KEYINPUT87), .A3(new_n381_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n283_), .B1(new_n338_), .B2(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n283_), .B2(KEYINPUT90), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  OAI221_X1 g189(.A(new_n283_), .B1(KEYINPUT90), .B2(new_n388_), .C1(new_n338_), .C2(new_n386_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(KEYINPUT93), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n392_), .B(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n338_), .A2(new_n386_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n397_), .A2(KEYINPUT28), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(KEYINPUT28), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G22gat), .B(G50gat), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n396_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT94), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n396_), .A2(KEYINPUT94), .A3(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n393_), .B1(new_n392_), .B2(KEYINPUT92), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n409_), .B1(KEYINPUT92), .B2(new_n392_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n392_), .A2(KEYINPUT92), .A3(new_n393_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n410_), .B(new_n411_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n384_), .A2(new_n385_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n408_), .A2(new_n382_), .A3(new_n412_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n316_), .B(new_n359_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n384_), .A2(new_n385_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n408_), .A2(new_n412_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  OR3_X1    g218(.A1(new_n352_), .A2(new_n419_), .A3(new_n357_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n342_), .A2(new_n347_), .A3(new_n318_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n357_), .B(new_n421_), .C1(new_n351_), .C2(new_n318_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n352_), .B2(new_n357_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n306_), .A2(new_n307_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT97), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n306_), .A2(KEYINPUT97), .A3(new_n307_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n424_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n304_), .A2(KEYINPUT32), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n312_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n294_), .A2(new_n299_), .A3(new_n430_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n431_), .A2(new_n358_), .A3(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n416_), .B(new_n418_), .C1(new_n429_), .C2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n242_), .B1(new_n415_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT69), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT65), .B(G85gat), .ZN(new_n438_));
  INV_X1    g237(.A(G92gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G99gat), .A2(G106gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(KEYINPUT10), .B(G99gat), .Z(new_n448_));
  INV_X1    g247(.A(G106gat), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n442_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G85gat), .B(G92gat), .Z(new_n452_));
  INV_X1    g251(.A(KEYINPUT8), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT7), .ZN(new_n455_));
  INV_X1    g254(.A(G99gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n449_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT66), .B1(new_n459_), .B2(new_n447_), .ZN(new_n460_));
  AND3_X1   g259(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT66), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n457_), .A4(new_n458_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n454_), .A2(new_n460_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n443_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT67), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(KEYINPUT6), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n444_), .A2(KEYINPUT67), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n467_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n458_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n444_), .A2(KEYINPUT67), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n468_), .A2(KEYINPUT6), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n443_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n471_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n453_), .B1(new_n478_), .B2(new_n452_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n451_), .B1(new_n466_), .B2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(G71gat), .A2(G78gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(G71gat), .A2(G78gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(KEYINPUT11), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(new_n484_), .B2(KEYINPUT11), .ZN(new_n487_));
  INV_X1    g286(.A(G64gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(G57gat), .ZN(new_n489_));
  INV_X1    g288(.A(G57gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G64gat), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n489_), .A2(new_n491_), .A3(new_n486_), .A4(KEYINPUT11), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n485_), .B1(new_n487_), .B2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n489_), .A2(new_n491_), .A3(KEYINPUT11), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT68), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n491_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT11), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n496_), .A2(new_n499_), .A3(new_n483_), .A4(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n494_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n480_), .A2(new_n502_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n451_), .B(new_n501_), .C1(new_n466_), .C2(new_n479_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(KEYINPUT12), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT12), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n480_), .A2(new_n506_), .A3(new_n502_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G230gat), .A2(G233gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT64), .Z(new_n510_));
  AOI21_X1  g309(.A(new_n436_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n510_), .ZN(new_n512_));
  AOI211_X1 g311(.A(KEYINPUT69), .B(new_n512_), .C1(new_n505_), .C2(new_n507_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT70), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n477_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n443_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n452_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT8), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n454_), .A2(new_n460_), .A3(new_n465_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n501_), .B1(new_n521_), .B2(new_n451_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n504_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n512_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G120gat), .B(G148gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT5), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G176gat), .B(G204gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n514_), .A2(new_n515_), .A3(new_n524_), .A4(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n504_), .A2(KEYINPUT12), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(new_n522_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n507_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n510_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT69), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n508_), .A2(new_n436_), .A3(new_n510_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n535_), .A2(new_n524_), .A3(new_n536_), .A4(new_n529_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT70), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n530_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n514_), .A2(new_n524_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n528_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT13), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(KEYINPUT71), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n539_), .A2(new_n541_), .A3(new_n544_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n530_), .A2(new_n538_), .B1(new_n540_), .B2(new_n528_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT34), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n206_), .B(new_n451_), .C1(new_n466_), .C2(new_n479_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n208_), .A2(new_n209_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n521_), .B2(new_n451_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n553_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n480_), .A2(new_n210_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n553_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n555_), .A4(new_n554_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT74), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT74), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n565_), .A3(new_n562_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G134gat), .B(G162gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT36), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n564_), .A2(new_n566_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT37), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n570_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT72), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n559_), .A2(new_n562_), .A3(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(new_n574_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n571_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n577_), .B1(new_n579_), .B2(KEYINPUT73), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT73), .ZN(new_n581_));
  AOI211_X1 g380(.A(new_n581_), .B(new_n571_), .C1(new_n559_), .C2(new_n562_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT37), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n578_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G127gat), .B(G155gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT17), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT78), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n230_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n501_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT80), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n593_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n593_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n596_), .A2(new_n502_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n596_), .A2(new_n502_), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT80), .B(new_n600_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n592_), .A2(KEYINPUT17), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n599_), .A2(new_n603_), .B1(new_n597_), .B2(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n585_), .A2(new_n586_), .A3(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n435_), .A2(new_n548_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n608_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612_));
  INV_X1    g411(.A(new_n359_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n212_), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n611_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n573_), .A2(new_n577_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n605_), .B(new_n617_), .C1(new_n415_), .C2(new_n434_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n242_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n548_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n359_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n612_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n615_), .A2(new_n624_), .A3(new_n625_), .ZN(G1324gat));
  INV_X1    g425(.A(new_n316_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n609_), .A2(new_n610_), .A3(new_n211_), .A4(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n622_), .A2(new_n627_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(new_n630_), .A3(G8gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n629_), .B2(G8gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n628_), .B(new_n634_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1325gat));
  INV_X1    g437(.A(new_n416_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n366_), .B1(new_n622_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT41), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n607_), .A2(new_n366_), .A3(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1326gat));
  AOI21_X1  g442(.A(new_n215_), .B1(new_n622_), .B2(new_n417_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT42), .Z(new_n645_));
  NAND3_X1  g444(.A1(new_n607_), .A2(new_n215_), .A3(new_n417_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(G29gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n621_), .A2(new_n605_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n415_), .A2(new_n434_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n585_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n586_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n651_), .B1(new_n652_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n655_), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT43), .B(new_n657_), .C1(new_n415_), .C2(new_n434_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n650_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT44), .B(new_n650_), .C1(new_n656_), .C2(new_n658_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n613_), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n648_), .B1(new_n663_), .B2(KEYINPUT103), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n664_), .B1(KEYINPUT103), .B2(new_n663_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n548_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n605_), .A2(new_n617_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n435_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n648_), .A3(new_n613_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n665_), .A2(new_n671_), .ZN(G1328gat));
  NOR2_X1   g471(.A1(new_n316_), .A2(G36gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n435_), .A2(new_n668_), .A3(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(KEYINPUT45), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(KEYINPUT45), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677_));
  OAI22_X1  g476(.A1(new_n675_), .A2(new_n676_), .B1(new_n677_), .B2(KEYINPUT46), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n661_), .A2(new_n627_), .A3(new_n662_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(G36gat), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n677_), .A2(KEYINPUT46), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1329gat));
  NAND3_X1  g481(.A1(new_n661_), .A2(new_n382_), .A3(new_n662_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G43gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n670_), .A2(new_n363_), .A3(new_n639_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(KEYINPUT47), .A3(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1330gat));
  AND4_X1   g489(.A1(G50gat), .A2(new_n661_), .A3(new_n417_), .A4(new_n662_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G50gat), .B1(new_n670_), .B2(new_n417_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1331gat));
  NAND3_X1  g492(.A1(new_n618_), .A2(new_n242_), .A3(new_n666_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n694_), .A2(new_n490_), .A3(new_n359_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT106), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n652_), .A2(new_n242_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n606_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n548_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT105), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(new_n359_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n696_), .B1(new_n701_), .B2(new_n490_), .ZN(G1332gat));
  OAI21_X1  g501(.A(G64gat), .B1(new_n694_), .B2(new_n316_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT48), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n627_), .A2(new_n488_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n700_), .B2(new_n705_), .ZN(G1333gat));
  OAI21_X1  g505(.A(G71gat), .B1(new_n694_), .B2(new_n416_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT49), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT49), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n416_), .A2(G71gat), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n708_), .A2(new_n709_), .B1(new_n700_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT107), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713_));
  OAI221_X1 g512(.A(new_n713_), .B1(new_n700_), .B2(new_n710_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1334gat));
  OAI21_X1  g514(.A(G78gat), .B1(new_n694_), .B2(new_n418_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT50), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n418_), .A2(G78gat), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT108), .Z(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n700_), .B2(new_n719_), .ZN(G1335gat));
  OR2_X1    g519(.A1(new_n548_), .A2(new_n667_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n697_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n613_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n656_), .A2(new_n658_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n605_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n548_), .A2(new_n619_), .A3(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n359_), .A2(new_n438_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n725_), .B1(new_n729_), .B2(new_n730_), .ZN(G1336gat));
  NAND3_X1  g530(.A1(new_n724_), .A2(new_n439_), .A3(new_n627_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n729_), .A2(new_n627_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n439_), .ZN(G1337gat));
  AND2_X1   g533(.A1(new_n382_), .A2(new_n448_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n724_), .A2(new_n735_), .B1(new_n736_), .B2(KEYINPUT51), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n736_), .A2(KEYINPUT51), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n726_), .A2(new_n639_), .A3(new_n728_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G99gat), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n737_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n738_), .B1(new_n737_), .B2(new_n740_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1338gat));
  XNOR2_X1  g542(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n417_), .B(new_n728_), .C1(new_n656_), .C2(new_n658_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(G106gat), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n745_), .A3(G106gat), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n722_), .A2(new_n723_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n697_), .A2(KEYINPUT109), .A3(new_n721_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n449_), .B(new_n417_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n744_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n749_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n753_), .B(new_n744_), .C1(new_n755_), .C2(new_n747_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n754_), .A2(new_n757_), .ZN(G1339gat));
  INV_X1    g557(.A(KEYINPUT59), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n548_), .A2(new_n606_), .A3(new_n242_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n548_), .A2(new_n606_), .A3(KEYINPUT112), .A4(new_n242_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(KEYINPUT54), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n760_), .A2(new_n761_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n242_), .B1(new_n530_), .B2(new_n538_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n535_), .A2(new_n769_), .A3(new_n536_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n505_), .A2(new_n512_), .A3(new_n507_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT113), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n505_), .A2(new_n773_), .A3(new_n512_), .A4(new_n507_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n512_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n772_), .A2(new_n774_), .B1(KEYINPUT55), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n770_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n528_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n779_), .B(new_n529_), .C1(new_n770_), .C2(new_n776_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n768_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT114), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n768_), .B(new_n783_), .C1(new_n778_), .C2(new_n780_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n239_), .B1(new_n235_), .B2(new_n228_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n227_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n233_), .A2(new_n229_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT115), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n232_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n785_), .B(new_n791_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n546_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n782_), .A2(new_n784_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n616_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(KEYINPUT57), .A3(new_n616_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n793_), .B1(new_n538_), .B2(new_n530_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n800_), .B(KEYINPUT58), .C1(new_n778_), .C2(new_n780_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n655_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n778_), .A2(new_n780_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT58), .B1(new_n803_), .B2(new_n800_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n798_), .A2(new_n799_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n767_), .B1(new_n807_), .B2(new_n605_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n627_), .A2(new_n359_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n414_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n759_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n810_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n805_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n727_), .B1(new_n813_), .B2(new_n799_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT59), .B(new_n812_), .C1(new_n814_), .C2(new_n767_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n242_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(G113gat), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT116), .B(new_n812_), .C1(new_n814_), .C2(new_n767_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n619_), .A2(new_n817_), .ZN(new_n822_));
  OAI22_X1  g621(.A1(new_n816_), .A2(new_n817_), .B1(new_n821_), .B2(new_n822_), .ZN(G1340gat));
  INV_X1    g622(.A(G120gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n548_), .B2(KEYINPUT60), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n824_), .A2(KEYINPUT60), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n819_), .A2(new_n820_), .A3(new_n825_), .A4(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n548_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(new_n824_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT117), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n827_), .C1(new_n828_), .C2(new_n824_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1341gat));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n819_), .A2(new_n820_), .A3(new_n834_), .A4(new_n727_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n605_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n834_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT118), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(new_n835_), .C1(new_n836_), .C2(new_n834_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1342gat));
  AOI21_X1  g640(.A(new_n657_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n842_));
  INV_X1    g641(.A(G134gat), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n617_), .A2(new_n843_), .ZN(new_n844_));
  OAI22_X1  g643(.A1(new_n842_), .A2(new_n843_), .B1(new_n821_), .B2(new_n844_), .ZN(G1343gat));
  INV_X1    g644(.A(new_n413_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n809_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n808_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n619_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT119), .B(G141gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1344gat));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n666_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g652(.A1(new_n807_), .A2(new_n605_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n767_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n856_), .A2(new_n413_), .A3(new_n727_), .A4(new_n809_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT120), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n848_), .A2(new_n859_), .A3(new_n727_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n858_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1346gat));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n848_), .A2(new_n326_), .A3(new_n617_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n326_), .B1(new_n848_), .B2(new_n655_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n865_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n856_), .A2(new_n413_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n870_), .A2(new_n657_), .A3(new_n847_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT121), .B(new_n866_), .C1(new_n871_), .C2(new_n326_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n869_), .A2(new_n872_), .ZN(G1347gat));
  NOR2_X1   g672(.A1(new_n613_), .A2(new_n316_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n416_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n856_), .A2(new_n619_), .A3(new_n418_), .A4(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n258_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT122), .B1(new_n877_), .B2(G169gat), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n877_), .A2(G169gat), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT62), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n883_), .A2(new_n884_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n882_), .B1(new_n886_), .B2(new_n887_), .ZN(G1348gat));
  NAND4_X1  g687(.A1(new_n856_), .A2(new_n418_), .A3(new_n666_), .A4(new_n876_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n257_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n808_), .A2(new_n417_), .ZN(new_n893_));
  INV_X1    g692(.A(G176gat), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n893_), .A2(new_n894_), .A3(new_n666_), .A4(new_n876_), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n891_), .A2(new_n892_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n892_), .B1(new_n891_), .B2(new_n895_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1349gat));
  NAND2_X1  g697(.A1(new_n893_), .A2(new_n876_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n249_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n900_), .A2(new_n267_), .A3(new_n727_), .A4(new_n902_), .ZN(new_n903_));
  OAI22_X1  g702(.A1(new_n899_), .A2(new_n605_), .B1(new_n901_), .B2(G183gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n899_), .B2(new_n657_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n617_), .A2(new_n268_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n899_), .B2(new_n907_), .ZN(G1351gat));
  NOR2_X1   g707(.A1(new_n870_), .A2(new_n875_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n619_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n666_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n914_));
  INV_X1    g713(.A(G211gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n727_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT125), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n909_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n914_), .A2(new_n915_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1354gat));
  NOR2_X1   g719(.A1(new_n808_), .A2(new_n846_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n617_), .A3(new_n874_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n921_), .A2(KEYINPUT126), .A3(new_n617_), .A4(new_n874_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT127), .B(G218gat), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n657_), .A2(new_n927_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n926_), .A2(new_n927_), .B1(new_n909_), .B2(new_n928_), .ZN(G1355gat));
endmodule


