//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G211gat), .B(G218gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n203_), .A2(new_n204_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT91), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n214_), .B(KEYINPUT90), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT1), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT91), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n219_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT92), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n225_), .A2(new_n226_), .B1(new_n217_), .B2(new_n216_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n219_), .A2(new_n223_), .A3(KEYINPUT92), .A4(new_n224_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n213_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n211_), .A2(KEYINPUT3), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n211_), .A2(KEYINPUT3), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n212_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n230_), .A2(new_n231_), .A3(new_n233_), .A4(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(new_n220_), .A3(new_n224_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n229_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n210_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(G228gat), .A3(G233gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n242_), .B(new_n210_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n202_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n243_), .A3(new_n202_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n238_), .A2(new_n239_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT28), .B(G22gat), .ZN(new_n249_));
  INV_X1    g048(.A(G50gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n248_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT93), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n252_), .B1(new_n244_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n245_), .A2(new_n253_), .A3(new_n246_), .A4(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259_));
  INV_X1    g058(.A(G92gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT18), .B(G64gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT19), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT94), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT87), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT23), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n268_), .A2(KEYINPUT23), .ZN(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT86), .B(G183gat), .Z(new_n273_));
  OAI22_X1  g072(.A1(new_n271_), .A2(new_n272_), .B1(G190gat), .B2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT22), .B(G169gat), .ZN(new_n275_));
  INV_X1    g074(.A(G176gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT88), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n278_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT88), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n274_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G190gat), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n273_), .A2(KEYINPUT25), .ZN(new_n286_));
  NOR2_X1   g085(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n268_), .A2(new_n270_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT87), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n268_), .B(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n291_), .B2(new_n270_), .ZN(new_n292_));
  OR2_X1    g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n293_), .A2(KEYINPUT24), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT24), .A3(new_n278_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n288_), .A2(new_n292_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n284_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT20), .B1(new_n299_), .B2(new_n210_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n292_), .B1(G183gat), .B2(G190gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n279_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n272_), .B1(new_n291_), .B2(KEYINPUT23), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(new_n296_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT25), .B(G183gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT95), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n285_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(KEYINPUT96), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT96), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n310_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n302_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n267_), .A2(new_n300_), .B1(new_n312_), .B2(new_n210_), .ZN(new_n313_));
  OAI211_X1 g112(.A(KEYINPUT94), .B(KEYINPUT20), .C1(new_n299_), .C2(new_n210_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n266_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n210_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n316_), .B(new_n302_), .C1(new_n309_), .C2(new_n311_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT20), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n299_), .B2(new_n210_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n319_), .A3(new_n266_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT97), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n317_), .A2(new_n319_), .A3(KEYINPUT97), .A4(new_n266_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n263_), .B1(new_n315_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n300_), .A2(new_n267_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n312_), .A2(new_n210_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n314_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n265_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n263_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(new_n323_), .A4(new_n322_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n313_), .A2(new_n266_), .A3(new_n314_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n316_), .A2(new_n302_), .A3(new_n308_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n319_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n265_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(KEYINPUT27), .B(new_n331_), .C1(new_n339_), .C2(new_n330_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n299_), .B(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G71gat), .B(G99gat), .Z(new_n344_));
  XOR2_X1   g143(.A(KEYINPUT30), .B(G15gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n343_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G127gat), .B(G134gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351_));
  INV_X1    g150(.A(G43gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n350_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n347_), .B(new_n354_), .Z(new_n355_));
  NOR3_X1   g154(.A1(new_n258_), .A2(new_n341_), .A3(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G57gat), .B(G85gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n350_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n229_), .B2(new_n237_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n224_), .B1(new_n218_), .B2(KEYINPUT91), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n221_), .A2(new_n222_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n226_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n216_), .A2(new_n217_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n228_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n212_), .A3(new_n211_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(new_n236_), .A3(new_n350_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n363_), .A2(new_n370_), .A3(KEYINPUT4), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n376_), .B(new_n362_), .C1(new_n229_), .C2(new_n237_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n373_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT99), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n374_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n375_), .A2(KEYINPUT99), .A3(new_n373_), .A4(new_n377_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n361_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n361_), .A3(new_n381_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n356_), .A2(new_n386_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n257_), .A2(new_n385_), .A3(new_n341_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n315_), .A2(new_n324_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(new_n389_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n380_), .A2(new_n361_), .A3(new_n381_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(new_n382_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT101), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n384_), .A2(KEYINPUT33), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n380_), .A2(new_n398_), .A3(new_n361_), .A4(new_n381_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n325_), .A2(KEYINPUT98), .A3(new_n331_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT98), .B1(new_n325_), .B2(new_n331_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n361_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n375_), .A2(new_n377_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n405_), .B2(new_n372_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n401_), .A2(new_n402_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(KEYINPUT101), .B(new_n392_), .C1(new_n393_), .C2(new_n382_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n396_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n388_), .B1(new_n410_), .B2(new_n257_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n355_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n387_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT37), .ZN(new_n414_));
  XOR2_X1   g213(.A(G43gat), .B(G50gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(G29gat), .B(G36gat), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n416_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT15), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT64), .B(G85gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n260_), .A2(KEYINPUT9), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G99gat), .A2(G106gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT6), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(G99gat), .A3(G106gat), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n422_), .A2(new_n423_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT9), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G85gat), .B(G92gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT10), .B(G99gat), .ZN(new_n431_));
  OAI221_X1 g230(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .C1(G106gat), .C2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT66), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n430_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT8), .ZN(new_n435_));
  INV_X1    g234(.A(G99gat), .ZN(new_n436_));
  INV_X1    g235(.A(G106gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(KEYINPUT65), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT7), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n425_), .A2(new_n427_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT7), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n441_), .A2(new_n436_), .A3(new_n437_), .A4(KEYINPUT65), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n434_), .A2(new_n435_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT65), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(G99gat), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n441_), .B1(new_n446_), .B2(new_n437_), .ZN(new_n447_));
  NOR4_X1   g246(.A1(new_n445_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT69), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT69), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n439_), .A2(new_n450_), .A3(new_n442_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT67), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT68), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n425_), .A2(new_n427_), .A3(new_n453_), .A4(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n455_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n440_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n449_), .A2(new_n451_), .A3(new_n456_), .A4(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n435_), .B1(new_n459_), .B2(new_n434_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n444_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AOI211_X1 g261(.A(KEYINPUT70), .B(new_n435_), .C1(new_n459_), .C2(new_n434_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n432_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT72), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT72), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n466_), .B(new_n432_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n421_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n419_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G232gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  OAI22_X1  g271(.A1(new_n464_), .A2(new_n469_), .B1(KEYINPUT35), .B2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(KEYINPUT35), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT35), .B(new_n472_), .C1(new_n468_), .C2(new_n473_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G134gat), .B(G162gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT77), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G190gat), .B(G218gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT36), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n483_), .B(KEYINPUT78), .Z(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n478_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n482_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(KEYINPUT36), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n476_), .A2(new_n488_), .A3(new_n477_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n414_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(KEYINPUT79), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n489_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT80), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n484_), .B1(new_n478_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n476_), .A2(KEYINPUT80), .A3(new_n477_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n493_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n490_), .B1(new_n497_), .B2(new_n414_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT79), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n492_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G127gat), .B(G155gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(G211gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT16), .B(G183gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT83), .B1(new_n505_), .B2(KEYINPUT17), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT81), .B(G15gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G1gat), .A2(G8gat), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n507_), .A2(G22gat), .B1(KEYINPUT14), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n509_), .B1(G22gat), .B2(new_n507_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G1gat), .B(G8gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT82), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n510_), .B(new_n512_), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n506_), .B(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G231gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G71gat), .B(G78gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(G57gat), .B(G64gat), .Z(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n519_), .B2(KEYINPUT11), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n520_), .B1(KEYINPUT11), .B2(new_n519_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n517_), .A3(KEYINPUT11), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n505_), .A2(KEYINPUT17), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n516_), .B2(new_n523_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n501_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(KEYINPUT12), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n467_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n451_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n450_), .B1(new_n439_), .B2(new_n442_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n434_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT8), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT70), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n460_), .A2(new_n461_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(new_n444_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n466_), .B1(new_n539_), .B2(new_n432_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n531_), .B1(new_n532_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT73), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n464_), .A2(new_n523_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT12), .B1(new_n464_), .B2(new_n523_), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n541_), .A2(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G230gat), .A2(G233gat), .ZN(new_n546_));
  AOI211_X1 g345(.A(new_n542_), .B(new_n530_), .C1(new_n465_), .C2(new_n467_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n546_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT71), .B1(new_n464_), .B2(new_n523_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n543_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n464_), .A2(KEYINPUT71), .A3(new_n523_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n550_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G176gat), .B(G204gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(G120gat), .B(G148gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n549_), .A2(new_n554_), .A3(new_n560_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT75), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n564_), .B1(new_n565_), .B2(KEYINPUT13), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n562_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n419_), .B(KEYINPUT84), .Z(new_n572_));
  INV_X1    g371(.A(new_n513_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT85), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(G229gat), .A3(G233gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n573_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n420_), .A2(new_n513_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G169gat), .B(G197gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n576_), .A2(new_n581_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n571_), .A2(new_n590_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n413_), .A2(new_n529_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(G1gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n385_), .B(KEYINPUT103), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT38), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT104), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n570_), .B2(new_n589_), .ZN(new_n599_));
  AOI211_X1 g398(.A(KEYINPUT104), .B(new_n590_), .C1(new_n566_), .C2(new_n569_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT105), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n497_), .B(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n527_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n599_), .A2(new_n600_), .A3(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n604_), .A2(new_n413_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n593_), .B1(new_n605_), .B2(new_n385_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n597_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n596_), .B2(new_n595_), .ZN(G1324gat));
  NOR2_X1   g407(.A1(new_n599_), .A2(new_n600_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n603_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n609_), .A2(new_n413_), .A3(new_n341_), .A4(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT106), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n604_), .A2(KEYINPUT106), .A3(new_n341_), .A4(new_n413_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .A4(G8gat), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT107), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n613_), .A2(G8gat), .A3(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT39), .ZN(new_n620_));
  INV_X1    g419(.A(G8gat), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n622_), .A2(KEYINPUT107), .A3(new_n614_), .A4(new_n615_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n618_), .A2(new_n620_), .A3(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n592_), .A2(new_n621_), .A3(new_n341_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  NAND2_X1  g428(.A1(new_n605_), .A2(new_n412_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G15gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT109), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT109), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n631_), .B(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT41), .ZN(new_n637_));
  INV_X1    g436(.A(G15gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n592_), .A2(new_n638_), .A3(new_n412_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT110), .Z(new_n640_));
  NAND3_X1  g439(.A1(new_n634_), .A2(new_n637_), .A3(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n605_), .B2(new_n258_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT42), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n592_), .A2(new_n642_), .A3(new_n258_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1327gat));
  NOR2_X1   g445(.A1(new_n602_), .A2(new_n527_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n413_), .A2(new_n591_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT111), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n413_), .A2(KEYINPUT111), .A3(new_n591_), .A4(new_n647_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G29gat), .B1(new_n652_), .B2(new_n385_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n609_), .A2(new_n528_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n413_), .B2(new_n501_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n413_), .A2(new_n655_), .A3(new_n501_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(KEYINPUT44), .ZN(new_n660_));
  INV_X1    g459(.A(G29gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n594_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(KEYINPUT44), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n653_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n650_), .A2(new_n666_), .A3(new_n341_), .A4(new_n651_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT45), .ZN(new_n668_));
  INV_X1    g467(.A(new_n341_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n654_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n658_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n656_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(new_n664_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT46), .B(new_n668_), .C1(new_n675_), .C2(new_n666_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n666_), .B1(new_n674_), .B2(new_n664_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n667_), .B(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n676_), .A2(new_n681_), .ZN(G1329gat));
  NAND2_X1  g481(.A1(new_n652_), .A2(new_n412_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n352_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n664_), .ZN(new_n685_));
  OAI211_X1 g484(.A(G43gat), .B(new_n412_), .C1(new_n659_), .C2(KEYINPUT44), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT47), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT47), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n684_), .B(new_n689_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1330gat));
  AOI21_X1  g490(.A(G50gat), .B1(new_n652_), .B2(new_n258_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n660_), .A2(new_n250_), .A3(new_n257_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n664_), .ZN(G1331gat));
  NOR2_X1   g493(.A1(new_n570_), .A2(new_n589_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n413_), .A2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(new_n529_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G57gat), .B1(new_n697_), .B2(new_n594_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT112), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n610_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT113), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n385_), .A2(G57gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(G1332gat));
  INV_X1    g502(.A(G64gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n697_), .A2(new_n704_), .A3(new_n341_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n701_), .A2(new_n341_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G64gat), .ZN(new_n708_));
  AOI211_X1 g507(.A(KEYINPUT48), .B(new_n704_), .C1(new_n701_), .C2(new_n341_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1333gat));
  INV_X1    g509(.A(G71gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n697_), .A2(new_n711_), .A3(new_n412_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT49), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n701_), .A2(new_n412_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(G71gat), .ZN(new_n715_));
  AOI211_X1 g514(.A(KEYINPUT49), .B(new_n711_), .C1(new_n701_), .C2(new_n412_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1334gat));
  INV_X1    g516(.A(G78gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n697_), .A2(new_n718_), .A3(new_n258_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n701_), .A2(new_n258_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(G78gat), .ZN(new_n722_));
  AOI211_X1 g521(.A(KEYINPUT50), .B(new_n718_), .C1(new_n701_), .C2(new_n258_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1335gat));
  NAND2_X1  g523(.A1(new_n696_), .A2(new_n647_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT114), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G85gat), .B1(new_n727_), .B2(new_n594_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n657_), .A2(new_n658_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n570_), .A2(new_n527_), .A3(new_n589_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n385_), .A2(new_n422_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n728_), .B1(new_n732_), .B2(new_n733_), .ZN(G1336gat));
  AOI21_X1  g533(.A(G92gat), .B1(new_n727_), .B2(new_n341_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n669_), .A2(new_n260_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n732_), .B2(new_n736_), .ZN(G1337gat));
  INV_X1    g536(.A(new_n431_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n727_), .A2(new_n738_), .A3(new_n412_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G99gat), .B1(new_n731_), .B2(new_n355_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n740_), .A3(new_n742_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1338gat));
  NOR2_X1   g545(.A1(new_n257_), .A2(G106gat), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n727_), .A2(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n258_), .B(new_n730_), .C1(new_n671_), .C2(new_n656_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(G106gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(G106gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT53), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n748_), .B(new_n755_), .C1(new_n752_), .C2(new_n751_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1339gat));
  NAND2_X1  g556(.A1(new_n575_), .A2(new_n580_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n579_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n758_), .B(new_n585_), .C1(new_n580_), .C2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(new_n588_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n563_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n544_), .A2(new_n543_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n530_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(KEYINPUT73), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n765_), .A2(new_n550_), .A3(new_n547_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n550_), .B1(new_n765_), .B2(new_n547_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(KEYINPUT55), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NOR4_X1   g568(.A1(new_n765_), .A2(new_n547_), .A3(new_n769_), .A4(new_n550_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n561_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n546_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n549_), .B1(new_n774_), .B2(new_n769_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n770_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n561_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n762_), .B1(new_n773_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT58), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n761_), .A2(new_n563_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n561_), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n772_), .B(new_n560_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(KEYINPUT116), .A3(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n781_), .A2(new_n787_), .A3(KEYINPUT117), .A4(new_n501_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n589_), .A2(new_n563_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n773_), .B2(new_n778_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n564_), .A2(new_n761_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n602_), .B(KEYINPUT57), .C1(new_n790_), .C2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n602_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n788_), .A2(new_n792_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n785_), .A2(KEYINPUT116), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n500_), .B1(new_n797_), .B2(KEYINPUT58), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT117), .B1(new_n798_), .B2(new_n787_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n528_), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n500_), .A2(new_n527_), .A3(new_n590_), .A4(new_n570_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT54), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n356_), .A2(new_n594_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n804_), .A2(KEYINPUT119), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n795_), .A2(new_n792_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n798_), .A2(new_n787_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n527_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n802_), .ZN(new_n814_));
  OAI221_X1 g613(.A(new_n810_), .B1(KEYINPUT119), .B2(new_n804_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(G113gat), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n590_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n807_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n806_), .B2(new_n590_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1340gat));
  NOR2_X1   g619(.A1(new_n570_), .A2(KEYINPUT60), .ZN(new_n821_));
  MUX2_X1   g620(.A(new_n821_), .B(KEYINPUT60), .S(G120gat), .Z(new_n822_));
  NAND3_X1  g621(.A1(new_n803_), .A2(new_n805_), .A3(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT120), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n804_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n815_), .B(new_n571_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G120gat), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n828_), .ZN(G1341gat));
  NAND2_X1  g628(.A1(new_n527_), .A2(G127gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT121), .Z(new_n831_));
  NAND3_X1  g630(.A1(new_n807_), .A2(new_n815_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(G127gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n806_), .B2(new_n528_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1342gat));
  INV_X1    g634(.A(G134gat), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n500_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n807_), .A2(new_n815_), .A3(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n806_), .B2(new_n602_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1343gat));
  AOI21_X1  g639(.A(new_n412_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n662_), .A2(new_n257_), .A3(new_n341_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n589_), .A3(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g643(.A1(new_n841_), .A2(new_n571_), .A3(new_n842_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g645(.A1(new_n841_), .A2(new_n527_), .A3(new_n842_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT61), .B(G155gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1346gat));
  INV_X1    g648(.A(new_n602_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n803_), .A2(new_n355_), .A3(new_n850_), .A4(new_n842_), .ZN(new_n851_));
  INV_X1    g650(.A(G162gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(KEYINPUT122), .A3(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n841_), .A2(G162gat), .A3(new_n501_), .A4(new_n842_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT122), .B1(new_n851_), .B2(new_n852_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1347gat));
  NOR4_X1   g656(.A1(new_n594_), .A2(new_n258_), .A3(new_n669_), .A4(new_n355_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G169gat), .B1(new_n859_), .B2(new_n590_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n859_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT124), .B(new_n858_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n865_), .A2(new_n275_), .A3(new_n589_), .A4(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(G169gat), .B(new_n861_), .C1(new_n859_), .C2(new_n590_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n863_), .A2(new_n867_), .A3(new_n868_), .ZN(G1348gat));
  NAND3_X1  g668(.A1(new_n865_), .A2(new_n571_), .A3(new_n866_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n803_), .A2(new_n858_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n570_), .A2(new_n276_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n870_), .A2(new_n276_), .B1(new_n871_), .B2(new_n872_), .ZN(G1349gat));
  AOI21_X1  g672(.A(new_n273_), .B1(new_n871_), .B2(new_n527_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n865_), .A2(new_n866_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n528_), .A2(new_n306_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(G1350gat));
  NAND3_X1  g676(.A1(new_n865_), .A2(new_n501_), .A3(new_n866_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G190gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n850_), .A2(new_n285_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT125), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n865_), .A2(new_n866_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1351gat));
  NOR3_X1   g682(.A1(new_n257_), .A2(new_n669_), .A3(new_n385_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n841_), .A2(new_n589_), .A3(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g685(.A1(new_n841_), .A2(new_n571_), .A3(new_n884_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g687(.A(new_n528_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n841_), .A2(new_n884_), .A3(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT126), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n890_), .B(new_n892_), .ZN(G1354gat));
  AND2_X1   g692(.A1(new_n841_), .A2(new_n884_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n850_), .ZN(new_n895_));
  INV_X1    g694(.A(G218gat), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n500_), .A2(new_n896_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n895_), .A2(new_n896_), .B1(new_n894_), .B2(new_n897_), .ZN(G1355gat));
endmodule


