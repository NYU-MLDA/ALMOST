//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OR2_X1    g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT24), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(KEYINPUT24), .A3(new_n206_), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n203_), .A2(new_n205_), .A3(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT26), .B(G190gat), .Z(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT22), .B(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n214_), .A2(new_n206_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT30), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G227gat), .A2(G233gat), .ZN(new_n221_));
  INV_X1    g020(.A(G15gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(G71gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(G99gat), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n225_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G127gat), .B(G134gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n226_), .A2(new_n231_), .A3(new_n227_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT79), .B(G43gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT31), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(new_n237_), .A3(new_n234_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G155gat), .A2(G162gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT80), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G155gat), .A2(G162gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(G141gat), .A2(G148gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT3), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n249_));
  INV_X1    g048(.A(G141gat), .ZN(new_n250_));
  INV_X1    g049(.A(G148gat), .ZN(new_n251_));
  OAI211_X1 g050(.A(KEYINPUT81), .B(new_n249_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n250_), .A2(new_n251_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT81), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT2), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n248_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT82), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n257_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n246_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n245_), .B(KEYINPUT1), .Z(new_n261_));
  AND2_X1   g060(.A1(new_n261_), .A2(new_n244_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n262_), .A2(new_n253_), .A3(new_n247_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT83), .B1(new_n260_), .B2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n256_), .A2(new_n257_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n256_), .A2(new_n257_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n244_), .B(new_n245_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT83), .ZN(new_n268_));
  INV_X1    g067(.A(new_n263_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n264_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT28), .B1(new_n271_), .B2(KEYINPUT29), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT84), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT29), .B1(new_n264_), .B2(new_n270_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n274_), .A2(new_n275_), .ZN(new_n278_));
  AOI211_X1 g077(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n264_), .C2(new_n270_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT84), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G22gat), .B(G50gat), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n277_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n264_), .A2(new_n270_), .A3(KEYINPUT29), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G197gat), .A2(G204gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT86), .B(G204gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(G197gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(G211gat), .B(G218gat), .Z(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT21), .A3(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT87), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n287_), .A2(G197gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT21), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(G197gat), .B2(G204gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n289_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(KEYINPUT21), .B2(new_n288_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G228gat), .A2(G233gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT29), .B1(new_n260_), .B2(new_n263_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n291_), .A2(new_n296_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n285_), .A2(new_n300_), .B1(new_n303_), .B2(new_n299_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NOR3_X1   g108(.A1(new_n283_), .A2(new_n284_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n285_), .A2(new_n300_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n303_), .A2(new_n299_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(new_n305_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT85), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n304_), .A2(new_n305_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n273_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n278_), .A2(new_n279_), .A3(KEYINPUT84), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n281_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n277_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n316_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n242_), .B1(new_n310_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n309_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n241_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT18), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n211_), .B(KEYINPUT89), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n210_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n208_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n218_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n332_), .B1(new_n297_), .B2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n302_), .A2(new_n219_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n338_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n302_), .A2(new_n219_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n332_), .B1(new_n302_), .B2(new_n336_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n341_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT90), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n343_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  AOI211_X1 g147(.A(KEYINPUT90), .B(new_n341_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n331_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n345_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n341_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT90), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n346_), .A2(new_n347_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n354_), .A2(new_n330_), .A3(new_n355_), .A4(new_n343_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT94), .B(KEYINPUT27), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n344_), .A2(new_n345_), .A3(new_n341_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n341_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT93), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  AOI211_X1 g162(.A(KEYINPUT93), .B(new_n341_), .C1(new_n338_), .C2(new_n342_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n331_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT27), .A3(new_n356_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n359_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n267_), .A2(new_n231_), .A3(new_n269_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT92), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n264_), .A2(new_n270_), .A3(new_n232_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT91), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT91), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n264_), .A2(new_n270_), .A3(new_n373_), .A4(new_n232_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n370_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n370_), .A2(new_n372_), .A3(KEYINPUT4), .A4(new_n374_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n264_), .A2(new_n270_), .A3(new_n379_), .A4(new_n232_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n376_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n377_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G85gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT0), .B(G57gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n377_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n367_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n354_), .A2(new_n355_), .A3(new_n343_), .A4(new_n394_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n377_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n388_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n399_), .A2(KEYINPUT33), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n377_), .A2(KEYINPUT33), .A3(new_n383_), .A4(new_n388_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n375_), .A2(new_n381_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n378_), .A2(new_n376_), .A3(new_n380_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(new_n389_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n403_), .A2(new_n406_), .A3(new_n356_), .A4(new_n350_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n401_), .B1(new_n402_), .B2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n242_), .B1(new_n324_), .B2(new_n323_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n326_), .A2(new_n393_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G1gat), .B(G8gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT75), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G15gat), .B(G22gat), .ZN(new_n413_));
  INV_X1    g212(.A(G1gat), .ZN(new_n414_));
  INV_X1    g213(.A(G8gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT14), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n411_), .A2(KEYINPUT75), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n411_), .A2(KEYINPUT75), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(new_n416_), .A3(new_n413_), .A4(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G43gat), .B(G50gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G36gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G29gat), .ZN(new_n426_));
  INV_X1    g225(.A(G29gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(G36gat), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n426_), .A2(new_n428_), .A3(KEYINPUT70), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT70), .B1(new_n426_), .B2(new_n428_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n424_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT70), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n427_), .A2(G36gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n425_), .A2(G29gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n426_), .A2(new_n428_), .A3(KEYINPUT70), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n423_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n431_), .A2(new_n437_), .A3(KEYINPUT15), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT15), .B1(new_n431_), .B2(new_n437_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n422_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G229gat), .A2(G233gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n431_), .A2(new_n437_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(new_n421_), .A3(new_n418_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n441_), .A2(KEYINPUT78), .A3(new_n442_), .A4(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n441_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n422_), .A2(new_n443_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n442_), .B1(new_n450_), .B2(new_n445_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G141gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G169gat), .B(G197gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  AND4_X1   g254(.A1(new_n446_), .A2(new_n449_), .A3(new_n452_), .A4(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n451_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n455_), .B1(new_n457_), .B2(new_n446_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT95), .B1(new_n410_), .B2(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n323_), .A2(new_n324_), .A3(new_n241_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n241_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n393_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n408_), .A2(new_n409_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT95), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n457_), .A2(new_n446_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n455_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n457_), .A2(new_n446_), .A3(new_n455_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n465_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n460_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G232gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT34), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT72), .B1(new_n475_), .B2(KEYINPUT35), .ZN(new_n476_));
  INV_X1    g275(.A(G106gat), .ZN(new_n477_));
  OR2_X1    g276(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT64), .ZN(new_n479_));
  NAND2_X1  g278(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n477_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n484_));
  INV_X1    g283(.A(G92gat), .ZN(new_n485_));
  OR2_X1    g284(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n484_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G99gat), .A2(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT6), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(G99gat), .A3(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n483_), .A2(new_n491_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n494_), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n492_), .A2(KEYINPUT6), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT66), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT66), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n493_), .A2(new_n495_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT7), .ZN(new_n504_));
  INV_X1    g303(.A(G99gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(new_n477_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n501_), .A2(new_n503_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G85gat), .B(G92gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n498_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  AOI211_X1 g311(.A(KEYINPUT8), .B(new_n510_), .C1(new_n508_), .C2(new_n496_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n497_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT15), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n443_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n438_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n476_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n508_), .A2(new_n496_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n498_), .A3(new_n511_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n502_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n506_), .A2(new_n507_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n510_), .B1(new_n523_), .B2(new_n503_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n520_), .B1(new_n524_), .B2(new_n498_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n525_), .A2(KEYINPUT71), .A3(new_n444_), .A4(new_n497_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n444_), .B(new_n497_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n518_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n475_), .A2(KEYINPUT35), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G134gat), .B(G162gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(KEYINPUT36), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n518_), .A2(new_n529_), .A3(new_n531_), .A4(new_n526_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT73), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n533_), .A2(new_n541_), .A3(new_n537_), .A4(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n533_), .A2(new_n538_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n536_), .B(KEYINPUT36), .Z(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n540_), .A2(new_n542_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(new_n544_), .A3(KEYINPUT37), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n556_));
  XOR2_X1   g355(.A(G71gat), .B(G78gat), .Z(new_n557_));
  OR2_X1    g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n557_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT76), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n561_), .B(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(new_n422_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n422_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G127gat), .B(G155gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT16), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G183gat), .B(G211gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n571_), .ZN(new_n573_));
  AND4_X1   g372(.A1(new_n565_), .A2(new_n566_), .A3(new_n572_), .A4(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n554_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n561_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n514_), .A2(new_n580_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n561_), .B(new_n497_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT12), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT12), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n514_), .A2(new_n584_), .A3(new_n580_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n579_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n578_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G120gat), .B(G148gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT5), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G176gat), .B(G204gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(KEYINPUT67), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n588_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n594_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n597_));
  XOR2_X1   g396(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT68), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n582_), .A2(KEYINPUT12), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n561_), .B1(new_n525_), .B2(new_n497_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n585_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n578_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n587_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n595_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n586_), .A2(new_n587_), .A3(new_n594_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n601_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n599_), .A2(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(KEYINPUT69), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(KEYINPUT69), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n577_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT77), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n473_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n414_), .A3(new_n392_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n410_), .A2(new_n551_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n611_), .A2(new_n471_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n576_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n392_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n618_), .A2(new_n619_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n620_), .A2(new_n627_), .A3(new_n628_), .ZN(G1324gat));
  NAND3_X1  g428(.A1(new_n617_), .A2(new_n415_), .A3(new_n367_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n621_), .A2(new_n367_), .A3(new_n624_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n631_), .A2(new_n632_), .A3(G8gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n631_), .B2(G8gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(G1325gat));
  OAI21_X1  g436(.A(G15gat), .B1(new_n625_), .B2(new_n241_), .ZN(new_n638_));
  XOR2_X1   g437(.A(KEYINPUT96), .B(KEYINPUT41), .Z(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT97), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n617_), .A2(new_n222_), .A3(new_n242_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(new_n640_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n641_), .A2(new_n642_), .A3(new_n643_), .ZN(G1326gat));
  NAND2_X1  g443(.A1(new_n323_), .A2(new_n324_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G22gat), .B1(new_n625_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT42), .ZN(new_n647_));
  INV_X1    g446(.A(G22gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n645_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n617_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(G1327gat));
  INV_X1    g450(.A(new_n551_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n576_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n611_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n473_), .A2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G29gat), .B1(new_n657_), .B2(new_n392_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n622_), .A2(new_n576_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n465_), .B2(new_n553_), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT43), .B(new_n554_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n659_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n410_), .B2(new_n554_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n465_), .A2(new_n660_), .A3(new_n553_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  AOI211_X1 g468(.A(new_n427_), .B(new_n626_), .C1(new_n669_), .C2(KEYINPUT44), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n658_), .B1(new_n665_), .B2(new_n670_), .ZN(G1328gat));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n672_), .A2(KEYINPUT98), .ZN(new_n673_));
  INV_X1    g472(.A(new_n367_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n669_), .B2(KEYINPUT44), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n425_), .B1(new_n675_), .B2(new_n665_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n674_), .A2(G36gat), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n410_), .A2(KEYINPUT95), .A3(new_n459_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n466_), .B1(new_n465_), .B2(new_n471_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n656_), .B(new_n677_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT45), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n473_), .A2(KEYINPUT45), .A3(new_n656_), .A4(new_n677_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n673_), .B1(new_n676_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n672_), .A2(KEYINPUT98), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT99), .Z(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n673_), .B(new_n687_), .C1(new_n676_), .C2(new_n684_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1329gat));
  NAND2_X1  g490(.A1(new_n669_), .A2(KEYINPUT44), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n665_), .A2(new_n692_), .A3(G43gat), .A4(new_n242_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n473_), .A2(new_n242_), .A3(new_n656_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n695_));
  INV_X1    g494(.A(G43gat), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n693_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT47), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n693_), .B(new_n701_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1330gat));
  INV_X1    g502(.A(G50gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n665_), .A2(new_n692_), .A3(new_n649_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(KEYINPUT101), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n706_), .B1(KEYINPUT101), .B2(new_n705_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n657_), .A2(new_n704_), .A3(new_n649_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1331gat));
  NAND4_X1  g508(.A1(new_n621_), .A2(new_n459_), .A3(new_n576_), .A4(new_n614_), .ZN(new_n710_));
  INV_X1    g509(.A(G57gat), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n626_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n410_), .A2(new_n471_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n577_), .A2(new_n611_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT102), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n626_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n717_), .B2(new_n716_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n712_), .B1(new_n719_), .B2(new_n711_), .ZN(G1332gat));
  OAI21_X1  g519(.A(G64gat), .B1(new_n710_), .B2(new_n674_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT48), .ZN(new_n722_));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n716_), .A2(new_n723_), .A3(new_n367_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1333gat));
  INV_X1    g524(.A(G71gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n716_), .A2(new_n726_), .A3(new_n242_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G71gat), .B1(new_n710_), .B2(new_n241_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(KEYINPUT49), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(KEYINPUT49), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT104), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n727_), .B(new_n733_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1334gat));
  OAI21_X1  g534(.A(G78gat), .B1(new_n710_), .B2(new_n645_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT50), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n645_), .A2(G78gat), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT105), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n716_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(G1335gat));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n742_));
  INV_X1    g541(.A(new_n614_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n654_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n713_), .A2(new_n742_), .A3(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n465_), .A2(new_n744_), .A3(new_n459_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT106), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n392_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n749_), .A2(KEYINPUT107), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(KEYINPUT107), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n611_), .A2(new_n471_), .A3(new_n576_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT108), .Z(new_n755_));
  AOI21_X1  g554(.A(new_n626_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n750_), .A2(new_n751_), .B1(new_n755_), .B2(new_n756_), .ZN(G1336gat));
  NAND3_X1  g556(.A1(new_n748_), .A2(new_n485_), .A3(new_n367_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n755_), .A2(new_n367_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(new_n485_), .ZN(G1337gat));
  OR2_X1    g559(.A1(new_n481_), .A2(new_n482_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n242_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n754_), .A2(new_n242_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n764_), .B(new_n765_), .C1(new_n766_), .C2(new_n505_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n505_), .B1(new_n754_), .B2(new_n242_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT110), .B1(new_n768_), .B2(new_n763_), .ZN(new_n769_));
  AND2_X1   g568(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n767_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n748_), .A2(new_n477_), .A3(new_n649_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n754_), .A2(new_n649_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(G106gat), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT52), .B(new_n477_), .C1(new_n754_), .C2(new_n649_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n774_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n450_), .A2(new_n445_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n455_), .B1(new_n786_), .B2(new_n442_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n441_), .A2(new_n445_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n442_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n470_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n606_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n586_), .A2(KEYINPUT55), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n583_), .A2(new_n579_), .A3(new_n585_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT114), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n583_), .A2(new_n797_), .A3(new_n579_), .A4(new_n585_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n793_), .A2(new_n794_), .A3(new_n796_), .A4(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n592_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n592_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n586_), .A2(new_n587_), .A3(new_n592_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n459_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n806_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n471_), .A2(new_n808_), .A3(KEYINPUT113), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n791_), .B1(new_n804_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n785_), .B1(new_n811_), .B2(new_n551_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n807_), .A2(new_n809_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT57), .B(new_n652_), .C1(new_n814_), .C2(new_n791_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n802_), .A2(KEYINPUT115), .A3(new_n803_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n470_), .A2(new_n789_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n808_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n592_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n817_), .A2(KEYINPUT58), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT58), .B1(new_n817_), .B2(new_n822_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n554_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n623_), .B1(new_n816_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n459_), .A2(new_n576_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n599_), .B2(new_n610_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n550_), .A2(new_n552_), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n832_));
  NAND4_X1  g631(.A1(new_n550_), .A2(new_n828_), .A3(KEYINPUT112), .A4(new_n552_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n832_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n554_), .A2(KEYINPUT112), .A3(new_n828_), .A4(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n826_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n674_), .A2(new_n392_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n322_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT59), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n592_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n844_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n800_), .A2(new_n821_), .A3(new_n801_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n819_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n843_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n817_), .A2(KEYINPUT58), .A3(new_n822_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n553_), .A3(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n837_), .B1(new_n852_), .B2(new_n623_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854_));
  INV_X1    g653(.A(new_n841_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n784_), .B1(new_n842_), .B2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n839_), .A2(KEYINPUT59), .A3(new_n841_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(KEYINPUT116), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n857_), .A2(new_n471_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G113gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n839_), .A2(new_n841_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n459_), .A2(G113gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(G1340gat));
  AOI21_X1  g664(.A(new_n743_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n866_));
  INV_X1    g665(.A(G120gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n611_), .B2(KEYINPUT60), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(KEYINPUT60), .B2(new_n867_), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n866_), .A2(new_n867_), .B1(new_n863_), .B2(new_n869_), .ZN(G1341gat));
  INV_X1    g669(.A(G127gat), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n623_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n857_), .A2(new_n860_), .A3(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n863_), .B2(new_n623_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n873_), .A2(KEYINPUT117), .A3(new_n874_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1342gat));
  AND2_X1   g678(.A1(new_n857_), .A2(new_n860_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT118), .B(G134gat), .Z(new_n881_));
  NOR2_X1   g680(.A1(new_n554_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(G134gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n839_), .A2(new_n551_), .A3(new_n841_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n880_), .A2(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1343gat));
  INV_X1    g684(.A(new_n840_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n461_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n887_), .A2(KEYINPUT119), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(KEYINPUT119), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n853_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n471_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n614_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT120), .B(G148gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1345gat));
  NAND2_X1  g694(.A1(new_n890_), .A2(new_n576_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1346gat));
  INV_X1    g697(.A(new_n890_), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n899_), .A2(G162gat), .A3(new_n652_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G162gat), .B1(new_n899_), .B2(new_n554_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1347gat));
  NOR3_X1   g701(.A1(new_n322_), .A2(new_n674_), .A3(new_n392_), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n839_), .A2(new_n471_), .A3(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904_), .B2(KEYINPUT121), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n839_), .A2(new_n903_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n459_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  OAI22_X1  g709(.A1(new_n905_), .A2(new_n908_), .B1(KEYINPUT123), .B2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n904_), .A2(KEYINPUT121), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n907_), .B1(new_n906_), .B2(new_n459_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n910_), .A2(KEYINPUT123), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n912_), .A2(G169gat), .A3(new_n913_), .A4(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n910_), .A2(KEYINPUT123), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n911_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n904_), .A2(new_n215_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1348gat));
  AND2_X1   g718(.A1(new_n839_), .A2(new_n903_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(new_n216_), .A3(new_n655_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G176gat), .B1(new_n906_), .B2(new_n743_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1349gat));
  OR3_X1    g722(.A1(new_n906_), .A2(new_n333_), .A3(new_n623_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n906_), .A2(new_n623_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(G183gat), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n906_), .B2(new_n554_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT125), .Z(new_n930_));
  NAND3_X1  g729(.A1(new_n920_), .A2(new_n210_), .A3(new_n551_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1351gat));
  NOR3_X1   g731(.A1(new_n674_), .A2(new_n325_), .A3(new_n392_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n839_), .A2(new_n933_), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n934_), .A2(KEYINPUT126), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(KEYINPUT126), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(G197gat), .B1(new_n937_), .B2(new_n471_), .ZN(new_n938_));
  INV_X1    g737(.A(G197gat), .ZN(new_n939_));
  AOI211_X1 g738(.A(new_n939_), .B(new_n459_), .C1(new_n935_), .C2(new_n936_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1352gat));
  AOI22_X1  g740(.A1(new_n937_), .A2(new_n614_), .B1(KEYINPUT127), .B2(G204gat), .ZN(new_n942_));
  INV_X1    g741(.A(G204gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n287_), .B1(KEYINPUT127), .B2(new_n943_), .ZN(new_n944_));
  AOI211_X1 g743(.A(new_n743_), .B(new_n944_), .C1(new_n935_), .C2(new_n936_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n942_), .A2(new_n945_), .ZN(G1353gat));
  OR2_X1    g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n947_), .B1(new_n937_), .B2(new_n576_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(KEYINPUT63), .B(G211gat), .ZN(new_n949_));
  AOI211_X1 g748(.A(new_n623_), .B(new_n949_), .C1(new_n935_), .C2(new_n936_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n948_), .A2(new_n950_), .ZN(G1354gat));
  INV_X1    g750(.A(G218gat), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n937_), .A2(new_n952_), .A3(new_n551_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n554_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n952_), .B2(new_n954_), .ZN(G1355gat));
endmodule


