//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT34), .ZN(new_n204_));
  XOR2_X1   g003(.A(G29gat), .B(G36gat), .Z(new_n205_));
  INV_X1    g004(.A(G43gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G29gat), .B(G36gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G43gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G50gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(G50gat), .A3(new_n209_), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n212_), .A2(KEYINPUT15), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT15), .B1(new_n212_), .B2(new_n213_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT64), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n218_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT9), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT10), .B(G99gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(G106gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n226_), .A2(KEYINPUT9), .ZN(new_n230_));
  OR3_X1    g029(.A1(new_n224_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT7), .ZN(new_n232_));
  INV_X1    g031(.A(G99gat), .ZN(new_n233_));
  INV_X1    g032(.A(G106gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .A4(KEYINPUT65), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236_));
  OAI22_X1  g035(.A1(new_n236_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n218_), .A2(new_n220_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n221_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n218_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n238_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n225_), .A2(new_n226_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n243_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n237_), .B(new_n235_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n244_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n245_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n231_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n224_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n246_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n248_), .A2(new_n249_), .A3(new_n245_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT69), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n216_), .B1(new_n253_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n213_), .ZN(new_n260_));
  AOI21_X1  g059(.A(G50gat), .B1(new_n207_), .B2(new_n209_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n251_), .A2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT35), .B(new_n204_), .C1(new_n259_), .C2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n214_), .A2(new_n215_), .ZN(new_n266_));
  AOI211_X1 g065(.A(new_n252_), .B(new_n254_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n255_), .A2(new_n256_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT69), .B1(new_n268_), .B2(new_n231_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n266_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n272_));
  INV_X1    g071(.A(new_n264_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .A4(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n265_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G162gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G190gat), .B(G218gat), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n277_), .A2(KEYINPUT71), .ZN(new_n278_));
  INV_X1    g077(.A(G134gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(KEYINPUT71), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n276_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(G162gat), .A3(new_n281_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT36), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT36), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(new_n286_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT73), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n275_), .A2(new_n292_), .A3(KEYINPUT74), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT74), .B1(new_n275_), .B2(new_n292_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n290_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n265_), .A2(new_n297_), .A3(new_n274_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n265_), .A2(new_n274_), .A3(KEYINPUT72), .A4(new_n297_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n202_), .B1(new_n296_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n275_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n265_), .A2(KEYINPUT75), .A3(new_n274_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n305_), .A2(new_n290_), .A3(new_n288_), .A4(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n307_), .A2(new_n202_), .A3(new_n302_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G127gat), .B(G155gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G183gat), .B(G211gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT17), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(KEYINPUT67), .A2(G57gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(KEYINPUT67), .A2(G57gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G64gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(G64gat), .A3(new_n318_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G71gat), .ZN(new_n324_));
  INV_X1    g123(.A(G78gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G71gat), .A2(G78gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n328_), .A2(KEYINPUT11), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(KEYINPUT11), .A3(new_n327_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n330_), .A2(KEYINPUT68), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(KEYINPUT68), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n323_), .A2(new_n329_), .A3(new_n331_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n332_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n321_), .B(new_n322_), .C1(KEYINPUT11), .C2(new_n328_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G231gat), .A2(G233gat), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n333_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT14), .ZN(new_n341_));
  AND2_X1   g140(.A1(KEYINPUT76), .A2(G8gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(KEYINPUT76), .A2(G8gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n344_), .B2(G1gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(G15gat), .B(G22gat), .Z(new_n346_));
  NOR3_X1   g145(.A1(new_n345_), .A2(KEYINPUT77), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT76), .B(G8gat), .ZN(new_n349_));
  INV_X1    g148(.A(G1gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT14), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n346_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n348_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(G1gat), .B1(new_n347_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT77), .B1(new_n345_), .B2(new_n346_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n348_), .A3(new_n352_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n350_), .A3(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(G8gat), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G8gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n357_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n350_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n359_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n340_), .A2(new_n358_), .A3(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n354_), .A2(G8gat), .A3(new_n357_), .ZN(new_n364_));
  AOI21_X1  g163(.A(G8gat), .B1(new_n354_), .B2(new_n357_), .ZN(new_n365_));
  OAI22_X1  g164(.A1(new_n364_), .A2(new_n365_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n316_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n314_), .A2(new_n315_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n363_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT79), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n363_), .A2(new_n371_), .A3(new_n366_), .A4(new_n368_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n367_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n309_), .A2(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(KEYINPUT80), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(KEYINPUT80), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT13), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n333_), .A2(new_n336_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT12), .B1(new_n251_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n251_), .A2(new_n381_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n381_), .A2(KEYINPUT12), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G230gat), .A2(G233gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n257_), .B(new_n381_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n388_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G120gat), .B(G148gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT5), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G176gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(G204gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n395_), .A2(KEYINPUT70), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n390_), .A2(new_n396_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n380_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n390_), .A2(new_n396_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(KEYINPUT13), .A3(new_n397_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n378_), .A2(new_n379_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G190gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT84), .B1(new_n405_), .B2(KEYINPUT26), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT25), .B(G183gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT26), .B(G190gat), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n406_), .B(new_n407_), .C1(new_n408_), .C2(KEYINPUT84), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(G169gat), .ZN(new_n412_));
  INV_X1    g211(.A(G176gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n409_), .A2(KEYINPUT85), .A3(new_n414_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT23), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(G183gat), .A3(G190gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT86), .ZN(new_n423_));
  INV_X1    g222(.A(G183gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT23), .B1(new_n424_), .B2(new_n405_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n422_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(G183gat), .B2(G190gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G169gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G197gat), .B(G204gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT21), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G211gat), .B(G218gat), .Z(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT91), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n440_), .A3(new_n437_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n436_), .A2(new_n437_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n434_), .A2(new_n435_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT20), .B1(new_n433_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT94), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n426_), .B1(G183gat), .B2(G190gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n431_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n408_), .A2(new_n407_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n451_), .A2(new_n414_), .A3(KEYINPUT95), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT95), .B1(new_n451_), .B2(new_n414_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n428_), .B(new_n419_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n446_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT19), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT94), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n460_), .B(KEYINPUT20), .C1(new_n433_), .C2(new_n446_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n448_), .A2(new_n456_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n433_), .A2(new_n446_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n455_), .A2(KEYINPUT101), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT101), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n442_), .B(new_n445_), .C1(new_n464_), .C2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(KEYINPUT100), .A2(KEYINPUT20), .ZN(new_n468_));
  OR2_X1    g267(.A1(KEYINPUT100), .A2(KEYINPUT20), .ZN(new_n469_));
  AND4_X1   g268(.A1(new_n463_), .A2(new_n467_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n462_), .B1(new_n470_), .B2(new_n459_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G8gat), .B(G36gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT18), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G64gat), .ZN(new_n474_));
  INV_X1    g273(.A(G92gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n471_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n463_), .ZN(new_n479_));
  OAI211_X1 g278(.A(KEYINPUT20), .B(new_n459_), .C1(new_n455_), .C2(new_n446_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n448_), .A2(new_n456_), .A3(new_n461_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n482_), .B2(new_n458_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n476_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n478_), .A2(KEYINPUT27), .A3(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G127gat), .B(G134gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(G113gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(G120gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT90), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G141gat), .A2(G148gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n490_), .B2(KEYINPUT89), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n491_), .A2(KEYINPUT3), .B1(new_n489_), .B2(new_n490_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G141gat), .A2(G148gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT2), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n492_), .B(new_n494_), .C1(KEYINPUT3), .C2(new_n491_), .ZN(new_n495_));
  INV_X1    g294(.A(G155gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n276_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT88), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G155gat), .A2(G162gat), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n499_), .B(KEYINPUT1), .Z(new_n502_));
  AOI21_X1  g301(.A(new_n490_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n493_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n488_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G120gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n487_), .B(new_n507_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n495_), .A2(new_n500_), .B1(new_n503_), .B2(new_n493_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(new_n510_), .A3(KEYINPUT4), .ZN(new_n511_));
  OR3_X1    g310(.A1(new_n508_), .A2(KEYINPUT4), .A3(new_n509_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G225gat), .A2(G233gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n511_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT96), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n506_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT96), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n511_), .A2(new_n512_), .A3(new_n518_), .A4(new_n514_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT98), .B(G1gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G85gat), .ZN(new_n524_));
  INV_X1    g323(.A(G29gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n523_), .B(new_n526_), .Z(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n520_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n516_), .A2(new_n527_), .A3(new_n517_), .A4(new_n519_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT27), .ZN(new_n533_));
  INV_X1    g332(.A(new_n484_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n483_), .A2(new_n476_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n485_), .A2(new_n532_), .A3(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G22gat), .B(G50gat), .Z(new_n538_));
  NOR3_X1   g337(.A1(new_n505_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT28), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT29), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n540_), .B1(new_n509_), .B2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n538_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT28), .B1(new_n505_), .B2(KEYINPUT29), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n509_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n538_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n446_), .B1(new_n509_), .B2(new_n541_), .ZN(new_n549_));
  INV_X1    g348(.A(G228gat), .ZN(new_n550_));
  INV_X1    g349(.A(G233gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  OAI221_X1 g352(.A(new_n446_), .B1(new_n550_), .B2(new_n551_), .C1(new_n509_), .C2(new_n541_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT93), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT93), .B1(new_n553_), .B2(new_n554_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n548_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT93), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(new_n543_), .A3(new_n547_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G78gat), .B(G106gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT92), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G15gat), .B(G43gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G227gat), .A2(G233gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  XOR2_X1   g365(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n567_));
  AND2_X1   g366(.A1(new_n433_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n433_), .A2(new_n567_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n566_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n433_), .A2(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n433_), .A2(new_n567_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n566_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G71gat), .B(G99gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT30), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n508_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n575_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n562_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n557_), .A2(new_n581_), .A3(new_n559_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n563_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n575_), .B(new_n578_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n557_), .A2(new_n581_), .A3(new_n559_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n581_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n476_), .A2(KEYINPUT32), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n529_), .A2(new_n530_), .B1(new_n483_), .B2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n471_), .A2(KEYINPUT32), .A3(new_n476_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n483_), .A2(new_n476_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n506_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n528_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n595_), .A2(KEYINPUT99), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(KEYINPUT99), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n593_), .A2(new_n599_), .A3(new_n484_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n530_), .B(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n592_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n585_), .A2(new_n586_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(new_n584_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n537_), .A2(new_n588_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n263_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT82), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n362_), .A2(new_n358_), .A3(new_n262_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT82), .B(new_n263_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n610_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n266_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n611_), .A3(new_n609_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G113gat), .B(G141gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT83), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n412_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(G197gat), .Z(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n614_), .A2(new_n616_), .A3(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n606_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n376_), .A2(new_n403_), .A3(new_n377_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT81), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n404_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n404_), .A2(KEYINPUT102), .A3(new_n627_), .A4(new_n629_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n632_), .A2(new_n350_), .A3(new_n531_), .A4(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n400_), .A2(new_n402_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n606_), .A2(new_n637_), .A3(new_n626_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n307_), .A2(new_n302_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n374_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n532_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n634_), .A2(new_n635_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n636_), .A2(new_n643_), .A3(new_n644_), .ZN(G1324gat));
  AND2_X1   g444(.A1(new_n485_), .A2(new_n536_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n632_), .A2(new_n349_), .A3(new_n647_), .A4(new_n633_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n649_));
  OAI211_X1 g448(.A(G8gat), .B(new_n649_), .C1(new_n642_), .C2(new_n646_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n648_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n648_), .A2(new_n653_), .A3(KEYINPUT40), .A4(new_n652_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1325gat));
  AND2_X1   g457(.A1(new_n632_), .A2(new_n633_), .ZN(new_n659_));
  INV_X1    g458(.A(G15gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n660_), .A3(new_n584_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G15gat), .B1(new_n642_), .B2(new_n580_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(new_n604_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(G22gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT105), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n659_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G22gat), .B1(new_n642_), .B2(new_n666_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT42), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n639_), .A2(new_n373_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n638_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n525_), .A3(new_n531_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n637_), .A2(new_n373_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n588_), .A2(new_n532_), .A3(new_n485_), .A4(new_n536_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n593_), .A2(new_n484_), .A3(new_n599_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n530_), .B(KEYINPUT33), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n679_), .A2(new_n680_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n605_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n309_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(new_n309_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n625_), .B(new_n677_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n275_), .A2(new_n292_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT74), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n302_), .A2(new_n692_), .A3(new_n293_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT37), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n307_), .A2(new_n202_), .A3(new_n302_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n606_), .B2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n683_), .A2(new_n684_), .A3(new_n309_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n699_), .A2(KEYINPUT44), .A3(new_n625_), .A4(new_n677_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n689_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n531_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n702_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT106), .B1(new_n702_), .B2(G29gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n676_), .B1(new_n703_), .B2(new_n704_), .ZN(G1328gat));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n689_), .A2(new_n700_), .A3(new_n647_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n689_), .A2(new_n700_), .A3(KEYINPUT107), .A4(new_n647_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(G36gat), .A3(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n674_), .A2(G36gat), .A3(new_n646_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT45), .Z(new_n713_));
  AOI211_X1 g512(.A(KEYINPUT108), .B(new_n706_), .C1(new_n711_), .C2(new_n713_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n716_));
  AND4_X1   g515(.A1(new_n715_), .A2(new_n711_), .A3(new_n716_), .A4(new_n713_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n714_), .A2(new_n717_), .ZN(G1329gat));
  AOI21_X1  g517(.A(G43gat), .B1(new_n675_), .B2(new_n584_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n580_), .A2(new_n206_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n701_), .B2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g521(.A1(new_n675_), .A2(new_n211_), .A3(new_n604_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n701_), .A2(new_n604_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n211_), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n403_), .A2(new_n625_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n606_), .A2(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n378_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n531_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n728_), .A2(new_n641_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n531_), .A2(G57gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(G1332gat));
  AOI21_X1  g532(.A(new_n320_), .B1(new_n731_), .B2(new_n647_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT48), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n729_), .A2(new_n320_), .A3(new_n647_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1333gat));
  AOI21_X1  g536(.A(new_n324_), .B1(new_n731_), .B2(new_n584_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT109), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT49), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n729_), .A2(new_n324_), .A3(new_n584_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1334gat));
  AOI21_X1  g541(.A(new_n325_), .B1(new_n731_), .B2(new_n604_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT50), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n729_), .A2(new_n325_), .A3(new_n604_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1335gat));
  AND2_X1   g545(.A1(new_n728_), .A2(new_n673_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n531_), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n373_), .B(new_n727_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n531_), .A2(G85gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT110), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n749_), .B2(new_n751_), .ZN(G1336gat));
  AOI21_X1  g551(.A(G92gat), .B1(new_n747_), .B2(new_n647_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n646_), .A2(new_n475_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n749_), .B2(new_n754_), .ZN(G1337gat));
  AOI21_X1  g554(.A(new_n233_), .B1(new_n749_), .B2(new_n584_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n580_), .A2(new_n228_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n747_), .B2(new_n757_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g558(.A1(new_n747_), .A2(new_n234_), .A3(new_n604_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n749_), .A2(new_n604_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(G106gat), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT52), .B(new_n234_), .C1(new_n749_), .C2(new_n604_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g565(.A1(new_n623_), .A2(new_n373_), .A3(new_n624_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n623_), .A2(KEYINPUT111), .A3(new_n373_), .A4(new_n624_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n403_), .C1(new_n303_), .C2(new_n308_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT54), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT113), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n775_), .A3(KEYINPUT54), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT112), .B1(new_n772_), .B2(KEYINPUT54), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n637_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .A4(new_n771_), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n774_), .A2(new_n776_), .B1(new_n777_), .B2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n387_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n388_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n384_), .A2(new_n386_), .A3(KEYINPUT55), .A4(new_n387_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n395_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT56), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n390_), .A2(new_n395_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n793_), .A3(new_n395_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n610_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n615_), .A2(new_n612_), .A3(new_n609_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n622_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n624_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n624_), .B2(new_n798_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n784_), .B1(new_n795_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n793_), .B1(new_n789_), .B2(new_n395_), .ZN(new_n805_));
  AOI211_X1 g604(.A(KEYINPUT56), .B(new_n394_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n624_), .A2(new_n798_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT114), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n800_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n807_), .A2(new_n810_), .A3(new_n792_), .A4(new_n783_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n804_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n309_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT116), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n791_), .A2(new_n625_), .A3(new_n792_), .A4(new_n794_), .ZN(new_n815_));
  OAI22_X1  g614(.A1(new_n801_), .A2(new_n802_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT57), .B1(new_n817_), .B2(new_n639_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n819_), .B(new_n640_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n812_), .A2(new_n822_), .A3(new_n309_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n814_), .A2(new_n821_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n782_), .B1(new_n824_), .B2(new_n374_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n647_), .A2(new_n532_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(new_n584_), .A3(new_n666_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828_), .B2(new_n625_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT117), .ZN(new_n830_));
  INV_X1    g629(.A(new_n828_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n774_), .A2(new_n776_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n777_), .A2(new_n781_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n821_), .A2(new_n813_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n373_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n827_), .A2(KEYINPUT59), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n831_), .A2(KEYINPUT59), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n625_), .A2(G113gat), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT118), .Z(new_n840_));
  AOI21_X1  g639(.A(new_n830_), .B1(new_n838_), .B2(new_n840_), .ZN(G1340gat));
  NOR2_X1   g640(.A1(new_n403_), .A2(G120gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n828_), .B1(KEYINPUT60), .B2(new_n842_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n838_), .A2(new_n637_), .A3(new_n843_), .ZN(new_n844_));
  OAI22_X1  g643(.A1(new_n844_), .A2(new_n507_), .B1(KEYINPUT60), .B2(new_n843_), .ZN(G1341gat));
  AOI21_X1  g644(.A(G127gat), .B1(new_n828_), .B2(new_n373_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n373_), .A2(G127gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT119), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n838_), .B2(new_n848_), .ZN(G1342gat));
  AOI21_X1  g648(.A(G134gat), .B1(new_n828_), .B2(new_n640_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n696_), .A2(new_n279_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT120), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n838_), .B2(new_n852_), .ZN(G1343gat));
  INV_X1    g652(.A(new_n826_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n825_), .A2(new_n583_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n625_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n637_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g658(.A(new_n640_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT57), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n822_), .B1(new_n812_), .B2(new_n309_), .ZN(new_n862_));
  AOI211_X1 g661(.A(KEYINPUT116), .B(new_n696_), .C1(new_n804_), .C2(new_n811_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n834_), .B1(new_n864_), .B2(new_n373_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n583_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n865_), .A2(new_n373_), .A3(new_n866_), .A4(new_n826_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT121), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n824_), .A2(new_n374_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n583_), .B1(new_n870_), .B2(new_n834_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n373_), .A4(new_n826_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n868_), .A2(new_n869_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n869_), .B1(new_n868_), .B2(new_n873_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n496_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n872_), .B1(new_n855_), .B2(new_n373_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n862_), .A2(new_n863_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n373_), .B1(new_n878_), .B2(new_n821_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n866_), .B(new_n826_), .C1(new_n879_), .C2(new_n782_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n880_), .A2(KEYINPUT121), .A3(new_n374_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT61), .B1(new_n877_), .B2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n868_), .A2(new_n869_), .A3(new_n873_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(G155gat), .A3(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n876_), .A2(new_n884_), .ZN(G1346gat));
  AOI21_X1  g684(.A(G162gat), .B1(new_n855_), .B2(new_n640_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n880_), .A2(new_n276_), .A3(new_n696_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1347gat));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n646_), .A2(new_n531_), .A3(new_n580_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT122), .B1(new_n891_), .B2(new_n626_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n893_), .A3(new_n625_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n836_), .A2(new_n889_), .A3(new_n666_), .A4(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n373_), .B1(new_n821_), .B2(new_n813_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n895_), .B(new_n666_), .C1(new_n782_), .C2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT123), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n896_), .A2(new_n899_), .A3(new_n900_), .A4(G169gat), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n896_), .A2(new_n899_), .A3(G169gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT62), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n901_), .A2(new_n902_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n903_), .A2(new_n905_), .A3(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n891_), .A2(new_n626_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT22), .B(G169gat), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n836_), .A2(new_n666_), .A3(new_n908_), .A4(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n910_), .ZN(G1348gat));
  NAND3_X1  g710(.A1(new_n836_), .A2(new_n666_), .A3(new_n890_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G176gat), .B1(new_n913_), .B2(new_n637_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n865_), .A2(new_n666_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT125), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n916_), .A2(new_n890_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n403_), .A2(new_n413_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n914_), .B1(new_n917_), .B2(new_n918_), .ZN(G1349gat));
  NOR3_X1   g718(.A1(new_n912_), .A2(new_n374_), .A3(new_n407_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n916_), .A2(new_n373_), .A3(new_n890_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n424_), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n912_), .B2(new_n696_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n640_), .A2(new_n408_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(KEYINPUT126), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n923_), .B1(new_n912_), .B2(new_n925_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT127), .ZN(G1351gat));
  NOR4_X1   g726(.A1(new_n825_), .A2(new_n531_), .A3(new_n583_), .A4(new_n646_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n625_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n637_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g731(.A1(new_n928_), .A2(new_n373_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT63), .B(G211gat), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n933_), .B2(new_n936_), .ZN(G1354gat));
  AOI21_X1  g736(.A(G218gat), .B1(new_n928_), .B2(new_n640_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n309_), .A2(G218gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n928_), .B2(new_n939_), .ZN(G1355gat));
endmodule


