//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G134gat), .ZN(new_n203_));
  INV_X1    g002(.A(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT7), .ZN(new_n207_));
  INV_X1    g006(.A(G99gat), .ZN(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT67), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT8), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n216_), .A2(new_n220_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(new_n214_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT10), .B(G99gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT64), .B1(new_n226_), .B2(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n208_), .A2(KEYINPUT10), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n208_), .A2(KEYINPUT10), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n228_), .B(new_n209_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n225_), .B1(new_n227_), .B2(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n233_));
  NOR2_X1   g032(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n217_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT66), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n219_), .B1(new_n218_), .B2(KEYINPUT9), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n238_), .B(new_n217_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n222_), .A2(new_n224_), .B1(new_n232_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G36gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G29gat), .ZN(new_n246_));
  INV_X1    g045(.A(G29gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G36gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(G43gat), .A2(G50gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G43gat), .A2(G50gat), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n246_), .B(new_n248_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n244_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n242_), .A2(new_n243_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n256_), .B2(new_n251_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT35), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G232gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT34), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n241_), .A2(new_n258_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n222_), .A2(new_n224_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n232_), .A2(new_n240_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n256_), .A2(new_n253_), .A3(new_n251_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n254_), .B1(new_n244_), .B2(new_n252_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT15), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT15), .B1(new_n267_), .B2(new_n268_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n266_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n262_), .A2(new_n259_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n263_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT76), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n263_), .A2(new_n271_), .A3(KEYINPUT76), .A4(new_n273_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT75), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n271_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT15), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT15), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(KEYINPUT75), .A3(new_n266_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(new_n285_), .A3(new_n263_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n286_), .A2(new_n272_), .ZN(new_n287_));
  OAI211_X1 g086(.A(KEYINPUT78), .B(new_n206_), .C1(new_n278_), .C2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n276_), .A2(new_n277_), .B1(new_n286_), .B2(new_n272_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n206_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT36), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n293_), .A3(new_n205_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n288_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT37), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT13), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G230gat), .A2(G233gat), .ZN(new_n299_));
  AND2_X1   g098(.A1(G57gat), .A2(G64gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G57gat), .A2(G64gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT11), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT68), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n304_), .B(KEYINPUT11), .C1(new_n300_), .C2(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  OR3_X1    g105(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT11), .ZN(new_n307_));
  XOR2_X1   g106(.A(G71gat), .B(G78gat), .Z(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n303_), .A2(new_n307_), .A3(new_n308_), .A4(new_n305_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT12), .ZN(new_n314_));
  OAI22_X1  g113(.A1(new_n241_), .A2(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(new_n241_), .B2(new_n312_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n310_), .A2(new_n311_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n313_), .A2(new_n314_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n266_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  AND4_X1   g119(.A1(new_n299_), .A2(new_n315_), .A3(new_n317_), .A4(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n299_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n266_), .A2(new_n318_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n241_), .A2(new_n312_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G120gat), .B(G148gat), .Z(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT71), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT72), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G176gat), .B(G204gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n329_), .B(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n322_), .A2(new_n326_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n333_), .B1(new_n322_), .B2(new_n326_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n298_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(KEYINPUT13), .A3(new_n334_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n206_), .B(KEYINPUT77), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n294_), .B(KEYINPUT37), .C1(new_n290_), .C2(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n297_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G231gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n312_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G8gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT79), .B(G8gat), .ZN(new_n349_));
  INV_X1    g148(.A(G1gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT14), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G15gat), .B(G22gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n348_), .A2(new_n353_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n345_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n345_), .A2(new_n357_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT17), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n362_));
  INV_X1    g161(.A(G155gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G183gat), .B(G211gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n364_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT82), .B(G127gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n367_), .A2(new_n368_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n361_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n369_), .A3(KEYINPUT17), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n360_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n358_), .A2(new_n374_), .A3(new_n359_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n377_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n343_), .A2(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT84), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G113gat), .B(G141gat), .ZN(new_n385_));
  INV_X1    g184(.A(G169gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G197gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n356_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n267_), .A2(new_n268_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n354_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(new_n284_), .B2(new_n357_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G229gat), .A2(G233gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n258_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n392_), .B1(new_n391_), .B2(new_n354_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n394_), .A2(new_n395_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n398_), .A2(new_n399_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n390_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n401_), .A3(new_n390_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G183gat), .A2(G190gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT23), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT23), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(G183gat), .A3(G190gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  INV_X1    g212(.A(G176gat), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n411_), .A2(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT101), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n416_), .A2(KEYINPUT101), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT87), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n408_), .A2(new_n410_), .A3(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n409_), .A2(KEYINPUT87), .A3(G183gat), .A4(G190gat), .ZN(new_n422_));
  OR3_X1    g221(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT99), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT99), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n421_), .A2(new_n426_), .A3(new_n422_), .A4(new_n423_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT25), .B(G183gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT26), .B(G190gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n386_), .A2(new_n414_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(KEYINPUT24), .A3(new_n416_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n428_), .A2(KEYINPUT100), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT100), .B1(new_n428_), .B2(new_n434_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n419_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G197gat), .B(G204gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT21), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G211gat), .B(G218gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT97), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT97), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n441_), .A2(new_n444_), .ZN(new_n446_));
  OAI22_X1  g245(.A1(new_n445_), .A2(new_n446_), .B1(new_n439_), .B2(new_n438_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n406_), .B1(new_n437_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT88), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n421_), .A2(new_n412_), .A3(new_n422_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n413_), .A2(new_n452_), .A3(new_n414_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n414_), .B1(new_n452_), .B2(KEYINPUT22), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G169gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n431_), .A2(new_n411_), .A3(new_n433_), .A4(new_n423_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n450_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(new_n450_), .A3(new_n457_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n443_), .A2(new_n447_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n449_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G226gat), .A2(G233gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT19), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT98), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n465_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n461_), .A2(new_n419_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n428_), .A2(new_n434_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n460_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n448_), .B1(new_n472_), .B2(new_n458_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT105), .B(KEYINPUT20), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n471_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  OAI22_X1  g274(.A1(new_n463_), .A2(new_n467_), .B1(new_n468_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT18), .B(G64gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G92gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n463_), .A2(new_n467_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n469_), .B1(new_n436_), .B2(new_n435_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n484_), .A2(KEYINPUT20), .A3(new_n468_), .A4(new_n473_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n480_), .A3(new_n485_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n482_), .A2(KEYINPUT27), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n466_), .B1(new_n449_), .B2(new_n462_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n485_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n481_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT27), .B1(new_n486_), .B2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G225gat), .A2(G233gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(G127gat), .B(G134gat), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT91), .B(G113gat), .ZN(new_n496_));
  INV_X1    g295(.A(G120gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G113gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT91), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(G113gat), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n500_), .A2(new_n502_), .A3(new_n497_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n495_), .B1(new_n498_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n500_), .A2(new_n502_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G120gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n496_), .A2(new_n497_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n494_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G155gat), .A2(G162gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT94), .B1(new_n510_), .B2(KEYINPUT1), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT1), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(G155gat), .A4(G162gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(KEYINPUT1), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n363_), .A2(new_n204_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n511_), .A2(new_n514_), .A3(new_n515_), .A4(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G141gat), .ZN(new_n518_));
  INV_X1    g317(.A(G148gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G141gat), .A2(G148gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT93), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(G141gat), .A3(G148gat), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n517_), .A2(new_n520_), .A3(new_n522_), .A4(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT2), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n522_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n520_), .A2(KEYINPUT3), .ZN(new_n529_));
  OR3_X1    g328(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .A4(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(new_n510_), .A3(new_n516_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n509_), .B1(new_n525_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT4), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n493_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n509_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n525_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n509_), .A2(new_n532_), .A3(new_n525_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(KEYINPUT4), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(KEYINPUT102), .B1(new_n535_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n539_), .A3(new_n493_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n540_), .A3(KEYINPUT102), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT0), .B(G57gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G85gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(G1gat), .B(G29gat), .Z(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .A4(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n472_), .B2(new_n458_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n459_), .A2(KEYINPUT30), .A3(new_n460_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT90), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT31), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n555_), .A2(new_n556_), .A3(KEYINPUT90), .A4(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n536_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT90), .B1(new_n555_), .B2(new_n556_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G15gat), .B(G43gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G71gat), .B(G99gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G227gat), .A2(G233gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT89), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n567_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT92), .B1(new_n564_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n557_), .A2(new_n558_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT92), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n570_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n559_), .A2(new_n509_), .A3(new_n561_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n563_), .A2(new_n572_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n572_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n559_), .A2(new_n509_), .A3(new_n561_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n509_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n578_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n577_), .A2(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n537_), .A2(KEYINPUT29), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G78gat), .B(G106gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n537_), .A2(KEYINPUT29), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n448_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n587_), .B(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT96), .B(G233gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(G228gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(G22gat), .B(G50gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n587_), .B(new_n588_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n583_), .B(new_n584_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n591_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n595_), .B1(new_n591_), .B2(new_n598_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n553_), .B1(new_n582_), .B2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n599_), .A2(new_n600_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n577_), .A3(new_n581_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n492_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n483_), .A2(new_n485_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT104), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n476_), .A2(KEYINPUT32), .A3(new_n480_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT104), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n483_), .A2(new_n610_), .A3(new_n485_), .A4(new_n606_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n608_), .A2(new_n553_), .A3(new_n609_), .A4(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n544_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n541_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n543_), .A4(new_n551_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n552_), .A2(KEYINPUT33), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n540_), .B(new_n493_), .C1(KEYINPUT4), .C2(new_n538_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n538_), .A2(new_n539_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT103), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n549_), .B(new_n619_), .C1(new_n621_), .C2(new_n493_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n618_), .A2(new_n486_), .A3(new_n490_), .A4(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n612_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n582_), .A2(new_n601_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n605_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n383_), .A2(KEYINPUT84), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n384_), .A2(new_n405_), .A3(new_n627_), .A4(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n553_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n629_), .A2(G1gat), .A3(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT38), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n627_), .A2(new_n405_), .A3(new_n340_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n295_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n633_), .A2(new_n634_), .A3(new_n381_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n350_), .B1(new_n635_), .B2(new_n553_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT106), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n637_), .ZN(G1324gat));
  INV_X1    g437(.A(new_n492_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(new_n641_), .A3(G8gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n640_), .B2(G8gat), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n349_), .ZN(new_n644_));
  OAI22_X1  g443(.A1(new_n642_), .A2(new_n643_), .B1(new_n629_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(G1325gat));
  NAND2_X1  g446(.A1(new_n635_), .A2(new_n582_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G15gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT41), .ZN(new_n650_));
  INV_X1    g449(.A(new_n582_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n629_), .A2(G15gat), .A3(new_n651_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n650_), .A2(new_n652_), .ZN(G1326gat));
  XNOR2_X1  g452(.A(new_n603_), .B(KEYINPUT107), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n635_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G22gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT42), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n654_), .A2(G22gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n629_), .B2(new_n659_), .ZN(G1327gat));
  NAND3_X1  g459(.A1(new_n340_), .A2(new_n381_), .A3(new_n405_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n297_), .A2(new_n342_), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT43), .B(new_n663_), .C1(new_n605_), .C2(new_n626_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n297_), .A2(new_n342_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n627_), .B2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n662_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT44), .B(new_n662_), .C1(new_n664_), .C2(new_n667_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n670_), .A2(G29gat), .A3(new_n553_), .A4(new_n671_), .ZN(new_n672_));
  AOI211_X1 g471(.A(new_n295_), .B(new_n661_), .C1(new_n605_), .C2(new_n626_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n247_), .B1(new_n674_), .B2(new_n630_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n672_), .A2(new_n675_), .ZN(G1328gat));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(KEYINPUT109), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n677_), .A2(KEYINPUT109), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n670_), .A2(new_n639_), .A3(new_n671_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G36gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n295_), .B1(new_n605_), .B2(new_n626_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n245_), .A3(new_n662_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT108), .B1(new_n683_), .B2(new_n492_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n673_), .A2(new_n685_), .A3(new_n245_), .A4(new_n639_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n684_), .A2(new_n686_), .A3(KEYINPUT45), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT45), .B1(new_n684_), .B2(new_n686_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI211_X1 g488(.A(new_n678_), .B(new_n679_), .C1(new_n681_), .C2(new_n689_), .ZN(new_n690_));
  AND4_X1   g489(.A1(KEYINPUT109), .A2(new_n681_), .A3(new_n677_), .A4(new_n689_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1329gat));
  NAND4_X1  g491(.A1(new_n670_), .A2(G43gat), .A3(new_n582_), .A4(new_n671_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n674_), .A2(new_n651_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(G43gat), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g495(.A1(new_n670_), .A2(new_n601_), .A3(new_n671_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n697_), .A2(KEYINPUT110), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(KEYINPUT110), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(G50gat), .A3(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n654_), .A2(G50gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n674_), .B2(new_n701_), .ZN(G1331gat));
  INV_X1    g501(.A(new_n340_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n403_), .B(new_n404_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n627_), .A2(new_n703_), .A3(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(new_n666_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G57gat), .B1(new_n707_), .B2(new_n553_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n627_), .A2(new_n295_), .A3(new_n703_), .A4(new_n705_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n709_), .A2(new_n630_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(G57gat), .B2(new_n710_), .ZN(G1332gat));
  INV_X1    g510(.A(G64gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n707_), .A2(new_n712_), .A3(new_n639_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714_));
  INV_X1    g513(.A(new_n709_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n639_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n716_), .B2(G64gat), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT48), .B(new_n712_), .C1(new_n715_), .C2(new_n639_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n713_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT111), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n709_), .B2(new_n651_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT49), .ZN(new_n722_));
  INV_X1    g521(.A(G71gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n707_), .A2(new_n723_), .A3(new_n582_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1334gat));
  INV_X1    g524(.A(G78gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n707_), .A2(new_n726_), .A3(new_n655_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G78gat), .B1(new_n709_), .B2(new_n654_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n728_), .A2(KEYINPUT112), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(KEYINPUT112), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(KEYINPUT50), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT50), .B1(new_n729_), .B2(new_n730_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT113), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n735_), .B(new_n727_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1335gat));
  NOR3_X1   g536(.A1(new_n340_), .A2(new_n382_), .A3(new_n405_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n682_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n553_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n664_), .A2(new_n667_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n738_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n630_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n741_), .B1(new_n744_), .B2(G85gat), .ZN(G1336gat));
  INV_X1    g544(.A(G92gat), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n743_), .A2(new_n746_), .A3(new_n492_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G92gat), .B1(new_n740_), .B2(new_n639_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1337gat));
  OAI21_X1  g548(.A(G99gat), .B1(new_n743_), .B2(new_n651_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n739_), .A2(new_n226_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(new_n651_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(KEYINPUT114), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n751_), .A2(new_n754_), .A3(new_n651_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n750_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g556(.A1(new_n740_), .A2(new_n209_), .A3(new_n601_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n601_), .B(new_n738_), .C1(new_n664_), .C2(new_n667_), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(G106gat), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n759_), .B2(G106gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  XOR2_X1   g562(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(G1339gat));
  AND2_X1   g564(.A1(new_n284_), .A2(new_n357_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT118), .B1(new_n766_), .B2(new_n393_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n394_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n395_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n396_), .A2(new_n397_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n395_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n389_), .A3(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(new_n404_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n315_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n323_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT55), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n322_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n776_), .A2(new_n780_), .A3(new_n323_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n333_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n321_), .B1(KEYINPUT55), .B2(new_n777_), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT56), .B(new_n784_), .C1(new_n786_), .C2(new_n781_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n334_), .B(new_n775_), .C1(new_n785_), .C2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n784_), .B1(new_n786_), .B2(new_n781_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n335_), .B1(new_n794_), .B2(new_n787_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n790_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n775_), .A3(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n791_), .A2(new_n666_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n394_), .A2(new_n395_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n398_), .A2(new_n399_), .ZN(new_n800_));
  AND4_X1   g599(.A1(new_n401_), .A2(new_n799_), .A3(new_n800_), .A4(new_n390_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n334_), .B1(new_n801_), .B2(new_n402_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n794_), .B2(new_n787_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n774_), .A2(new_n404_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n338_), .B2(new_n334_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n295_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT57), .B(new_n295_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n798_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n381_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n704_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n813_), .A2(new_n340_), .A3(new_n297_), .A4(new_n342_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n704_), .A2(new_n812_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817_));
  INV_X1    g616(.A(new_n815_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n343_), .A2(new_n817_), .A3(new_n818_), .A4(new_n813_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n811_), .A2(new_n820_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n639_), .A2(new_n630_), .A3(new_n651_), .ZN(new_n822_));
  XOR2_X1   g621(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n823_));
  NAND4_X1  g622(.A1(new_n821_), .A2(new_n603_), .A3(new_n822_), .A4(new_n823_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n810_), .A2(new_n381_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n822_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n825_), .A2(new_n601_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n824_), .B(new_n405_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G113gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n499_), .A3(new_n405_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT121), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(new_n834_), .A3(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1340gat));
  OAI211_X1 g635(.A(new_n824_), .B(new_n703_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G120gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n497_), .B1(new_n340_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n827_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n497_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT122), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n838_), .A2(new_n843_), .A3(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1341gat));
  NOR3_X1   g644(.A1(new_n825_), .A2(new_n601_), .A3(new_n381_), .ZN(new_n846_));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n822_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n827_), .A2(new_n828_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n849_), .A2(new_n382_), .A3(new_n824_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n850_), .B2(new_n847_), .ZN(G1342gat));
  AOI21_X1  g650(.A(G134gat), .B1(new_n827_), .B2(new_n634_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n849_), .A2(new_n666_), .A3(new_n824_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g653(.A1(new_n825_), .A2(new_n630_), .A3(new_n639_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n603_), .A2(new_n582_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n405_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(new_n518_), .ZN(G1344gat));
  NOR2_X1   g659(.A1(new_n857_), .A2(new_n340_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n519_), .ZN(G1345gat));
  NOR2_X1   g661(.A1(new_n857_), .A2(new_n381_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(new_n363_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n863_), .B(new_n865_), .ZN(G1346gat));
  NOR3_X1   g665(.A1(new_n857_), .A2(new_n204_), .A3(new_n663_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n855_), .A2(new_n634_), .A3(new_n856_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n204_), .B2(new_n868_), .ZN(G1347gat));
  NAND3_X1  g668(.A1(new_n639_), .A2(new_n630_), .A3(new_n582_), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n825_), .A2(new_n858_), .A3(new_n655_), .A4(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n413_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n871_), .B2(new_n386_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n874_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT124), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n873_), .A2(new_n879_), .A3(new_n876_), .A4(new_n874_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1348gat));
  NOR2_X1   g680(.A1(new_n870_), .A2(new_n340_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n821_), .A2(new_n414_), .A3(new_n654_), .A4(new_n882_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n821_), .A2(new_n603_), .A3(new_n882_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n414_), .ZN(G1349gat));
  INV_X1    g684(.A(new_n870_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G183gat), .B1(new_n846_), .B2(new_n886_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n825_), .A2(new_n655_), .A3(new_n870_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n381_), .A2(new_n429_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(G1350gat));
  NAND3_X1  g689(.A1(new_n888_), .A2(new_n634_), .A3(new_n430_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n888_), .A2(new_n666_), .ZN(new_n892_));
  INV_X1    g691(.A(G190gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(G1351gat));
  AOI21_X1  g693(.A(KEYINPUT125), .B1(new_n856_), .B2(new_n630_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n492_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n856_), .A2(KEYINPUT125), .A3(new_n630_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n821_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n858_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n388_), .ZN(G1352gat));
  INV_X1    g699(.A(new_n898_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n703_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n821_), .A2(new_n896_), .A3(new_n897_), .A4(new_n904_), .ZN(new_n905_));
  OR3_X1    g704(.A1(new_n905_), .A2(KEYINPUT126), .A3(new_n381_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT126), .B1(new_n905_), .B2(new_n381_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n906_), .A2(new_n910_), .A3(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1354gat));
  AOI21_X1  g711(.A(G218gat), .B1(new_n901_), .B2(new_n634_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n898_), .A2(new_n663_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(G218gat), .B2(new_n914_), .ZN(G1355gat));
endmodule


