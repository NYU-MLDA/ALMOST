//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G71gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G78gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n204_), .B2(KEYINPUT11), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n206_));
  INV_X1    g005(.A(G78gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n203_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n206_), .A2(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n205_), .B1(new_n211_), .B2(new_n202_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G231gat), .A2(G233gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n213_), .B(KEYINPUT74), .Z(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n212_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G1gat), .ZN(new_n217_));
  INV_X1    g016(.A(G8gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT72), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT72), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n222_), .B(KEYINPUT14), .C1(new_n217_), .C2(new_n218_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT73), .ZN(new_n225_));
  XOR2_X1   g024(.A(G1gat), .B(G8gat), .Z(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n224_), .A2(KEYINPUT73), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(KEYINPUT73), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n216_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT75), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G127gat), .B(G155gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G211gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT16), .B(G183gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n235_), .B(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(new_n240_), .A3(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT6), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n249_));
  OR3_X1    g048(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G85gat), .B(G92gat), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT8), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(KEYINPUT9), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT10), .B(G99gat), .Z(new_n257_));
  INV_X1    g056(.A(G106gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT9), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(G85gat), .A3(G92gat), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n256_), .A2(new_n259_), .A3(new_n261_), .A4(new_n248_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n251_), .A2(KEYINPUT8), .A3(new_n252_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n255_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n255_), .A2(KEYINPUT66), .A3(new_n262_), .A4(new_n263_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G29gat), .B(G36gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G43gat), .B(G50gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT15), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n246_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n264_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n271_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(KEYINPUT35), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n251_), .A2(KEYINPUT8), .A3(new_n252_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT8), .B1(new_n251_), .B2(new_n252_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT66), .B1(new_n280_), .B2(new_n262_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n267_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n272_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n283_), .A2(KEYINPUT69), .A3(KEYINPUT70), .A4(new_n275_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT34), .ZN(new_n285_));
  INV_X1    g084(.A(G232gat), .ZN(new_n286_));
  INV_X1    g085(.A(G233gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT34), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n273_), .A2(KEYINPUT69), .A3(new_n290_), .A4(new_n275_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n285_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n289_), .B1(new_n285_), .B2(new_n291_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n277_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n285_), .A2(new_n291_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n288_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n285_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(KEYINPUT35), .A3(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G190gat), .B(G218gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G134gat), .B(G162gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(KEYINPUT36), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n294_), .A2(new_n298_), .A3(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n301_), .B(KEYINPUT36), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT71), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n306_), .B1(new_n294_), .B2(new_n298_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT37), .B1(new_n304_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n294_), .A2(new_n298_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n305_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT37), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n294_), .A2(new_n298_), .A3(new_n303_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n245_), .B1(new_n308_), .B2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT76), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G230gat), .A2(G233gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n211_), .A2(new_n202_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n205_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n320_), .A2(new_n264_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n212_), .A2(new_n274_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n317_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT65), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n268_), .A2(KEYINPUT12), .A3(new_n320_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT12), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n212_), .B2(new_n274_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n212_), .A2(new_n274_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n329_), .A2(KEYINPUT67), .A3(new_n316_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT67), .B1(new_n329_), .B2(new_n316_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n324_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G120gat), .B(G148gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(G204gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(KEYINPUT5), .B(G176gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n333_), .B(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n339_));
  OR2_X1    g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(KEYINPUT68), .B2(KEYINPUT13), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n232_), .A2(new_n272_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n228_), .A2(new_n231_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n271_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT77), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G229gat), .A2(G233gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(KEYINPUT78), .Z(new_n349_));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n343_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n271_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n344_), .B(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n354_), .A2(new_n348_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT81), .B(G197gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT80), .B(G169gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G113gat), .B(G141gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n361_), .A2(KEYINPUT79), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n356_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n342_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT103), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT27), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G92gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT18), .B(G64gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G204gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(G197gat), .ZN(new_n372_));
  INV_X1    g171(.A(G197gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G204gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT21), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT21), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n372_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G211gat), .B(G218gat), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G197gat), .B(G204gat), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n381_), .A2(new_n379_), .A3(new_n377_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G169gat), .ZN(new_n384_));
  INV_X1    g183(.A(G176gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT22), .B(G169gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n387_), .B2(new_n385_), .ZN(new_n388_));
  INV_X1    g187(.A(G183gat), .ZN(new_n389_));
  INV_X1    g188(.A(G190gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT23), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(G183gat), .A3(G190gat), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n388_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT24), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT24), .B1(new_n384_), .B2(new_n385_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(new_n397_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n393_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n391_), .A2(new_n393_), .A3(new_n403_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT25), .B(G183gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT26), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G190gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n390_), .A2(KEYINPUT26), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n406_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n402_), .A2(new_n404_), .A3(new_n405_), .A4(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n383_), .A2(new_n396_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT91), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n382_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(KEYINPUT91), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n414_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n390_), .A2(KEYINPUT82), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G190gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n407_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n408_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n401_), .B1(new_n426_), .B2(KEYINPUT83), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT82), .B(G190gat), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n408_), .B(new_n406_), .C1(new_n428_), .C2(new_n407_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n394_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n404_), .B(new_n405_), .C1(G183gat), .C2(new_n428_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n427_), .A2(new_n431_), .B1(new_n432_), .B2(new_n388_), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT20), .B(new_n412_), .C1(new_n418_), .C2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT19), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n418_), .A2(new_n433_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n383_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n411_), .A2(new_n396_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n439_), .A2(new_n442_), .A3(KEYINPUT20), .A4(new_n436_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n370_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n434_), .A2(new_n436_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT100), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n439_), .A2(new_n442_), .A3(KEYINPUT20), .A4(new_n437_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n434_), .A2(KEYINPUT100), .A3(new_n436_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI211_X1 g249(.A(new_n366_), .B(new_n444_), .C1(new_n450_), .C2(new_n370_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n444_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n438_), .A2(new_n443_), .A3(new_n370_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT27), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n365_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n370_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(KEYINPUT27), .A3(new_n452_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n454_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(KEYINPUT103), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G78gat), .B(G106gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n461_), .B(KEYINPUT94), .Z(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G141gat), .A3(G148gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT2), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(KEYINPUT2), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n471_), .A2(new_n467_), .B1(G141gat), .B2(G148gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n466_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G155gat), .A2(G162gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT1), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G141gat), .A2(G148gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT85), .ZN(new_n480_));
  OR2_X1    g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT1), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n468_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT86), .B1(new_n483_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(G141gat), .A2(G148gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(KEYINPUT85), .B2(new_n479_), .ZN(new_n490_));
  INV_X1    g289(.A(G155gat), .ZN(new_n491_));
  INV_X1    g290(.A(G162gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n486_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n477_), .B1(new_n488_), .B2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n499_));
  AOI21_X1  g298(.A(new_n383_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT93), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G228gat), .A2(G233gat), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n496_), .B1(new_n495_), .B2(new_n486_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n487_), .A2(KEYINPUT86), .A3(new_n494_), .A4(new_n490_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n504_), .A2(new_n505_), .B1(new_n476_), .B2(new_n473_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n499_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n440_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n502_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT93), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n503_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512_));
  AOI221_X4 g311(.A(new_n512_), .B1(new_n473_), .B2(new_n476_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n504_), .A2(new_n505_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT88), .B1(new_n514_), .B2(new_n477_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT29), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n418_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n502_), .B(KEYINPUT90), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n462_), .B1(new_n511_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n501_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n508_), .A2(KEYINPUT93), .A3(new_n509_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n462_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n520_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n498_), .A2(new_n512_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n506_), .A2(KEYINPUT88), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT28), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G22gat), .B(G50gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n529_), .A2(new_n531_), .A3(new_n535_), .A4(new_n530_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n534_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n528_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(new_n536_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n534_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(KEYINPUT89), .A3(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n527_), .A2(new_n539_), .A3(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n537_), .A2(new_n538_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT95), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n526_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n461_), .B1(new_n511_), .B2(new_n519_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n523_), .A2(KEYINPUT95), .A3(new_n524_), .A4(new_n525_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n546_), .A2(new_n548_), .A3(new_n549_), .A4(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n545_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT96), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n545_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n433_), .B(KEYINPUT30), .ZN(new_n556_));
  XOR2_X1   g355(.A(G113gat), .B(G120gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(G127gat), .B(G134gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n560_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G15gat), .B(G43gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT31), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n561_), .A2(new_n562_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G71gat), .B(G99gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G227gat), .A2(G233gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n567_), .A2(new_n568_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n561_), .A2(new_n562_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n564_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n575_), .B2(new_n566_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n460_), .A2(new_n553_), .A3(new_n555_), .A4(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n573_), .A2(new_n576_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n451_), .A2(new_n454_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n545_), .A2(new_n554_), .A3(new_n551_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n554_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n579_), .B(new_n580_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT98), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n559_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n585_), .B1(new_n586_), .B2(KEYINPUT4), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n506_), .A2(new_n560_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(KEYINPUT4), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G225gat), .A2(G233gat), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT97), .Z(new_n591_));
  NAND2_X1  g390(.A1(new_n529_), .A2(new_n531_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT4), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n592_), .A2(KEYINPUT98), .A3(new_n593_), .A4(new_n559_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n587_), .A2(new_n589_), .A3(new_n591_), .A4(new_n594_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n595_), .A2(KEYINPUT99), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n586_), .A2(new_n588_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n590_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(KEYINPUT99), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G1gat), .B(G29gat), .ZN(new_n601_));
  INV_X1    g400(.A(G85gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT0), .B(G57gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n605_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .A4(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n606_), .A2(KEYINPUT102), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT102), .B1(new_n606_), .B2(new_n608_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n606_), .A2(new_n608_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n370_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n450_), .A2(KEYINPUT32), .A3(new_n613_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n438_), .A2(new_n443_), .B1(KEYINPUT32), .B2(new_n613_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT101), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(KEYINPUT101), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n612_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n608_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n595_), .B(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n624_), .A2(KEYINPUT33), .A3(new_n598_), .A4(new_n607_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n453_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n444_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .A4(new_n594_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n597_), .A2(new_n591_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n605_), .A3(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n622_), .A2(new_n625_), .A3(new_n627_), .A4(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n620_), .A2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n581_), .A2(new_n577_), .A3(new_n582_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n584_), .A2(new_n611_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n364_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n315_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n611_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n217_), .A3(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT38), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n310_), .A2(new_n312_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(new_n245_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n635_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n611_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n639_), .A2(new_n644_), .ZN(G1324gat));
  INV_X1    g444(.A(new_n643_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n460_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n218_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n636_), .A2(new_n218_), .A3(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n643_), .B2(new_n579_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT41), .Z(new_n655_));
  INV_X1    g454(.A(G15gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n636_), .A2(new_n656_), .A3(new_n577_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n581_), .A2(new_n582_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G22gat), .B1(new_n643_), .B2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  INV_X1    g461(.A(new_n659_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n636_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(G1327gat));
  NOR2_X1   g464(.A1(new_n634_), .A2(new_n640_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n342_), .A2(new_n363_), .A3(new_n245_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n637_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n308_), .A2(new_n313_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n584_), .A2(new_n611_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n632_), .A2(new_n633_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n677_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT105), .B(KEYINPUT43), .C1(new_n634_), .C2(new_n673_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n667_), .B(KEYINPUT104), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n683_), .A2(new_n684_), .A3(KEYINPUT44), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n611_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n671_), .B1(new_n689_), .B2(G29gat), .ZN(G1328gat));
  NOR2_X1   g489(.A1(new_n669_), .A2(G36gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n647_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT45), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n460_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n694_));
  INV_X1    g493(.A(G36gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT46), .B(new_n693_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  XNOR2_X1  g499(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT44), .B1(new_n683_), .B2(new_n684_), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT106), .B(new_n686_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n577_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G43gat), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n669_), .A2(G43gat), .A3(new_n579_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n701_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n701_), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n709_), .B(new_n706_), .C1(new_n704_), .C2(G43gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1330gat));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n663_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G50gat), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n669_), .A2(G50gat), .A3(new_n659_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n712_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT108), .B(new_n715_), .C1(new_n713_), .C2(G50gat), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1331gat));
  NOR2_X1   g518(.A1(new_n342_), .A2(new_n363_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n674_), .A2(new_n675_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n642_), .ZN(new_n722_));
  INV_X1    g521(.A(G57gat), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n611_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n315_), .A2(new_n721_), .A3(new_n720_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n637_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n726_), .B2(new_n723_), .ZN(G1332gat));
  OAI21_X1  g526(.A(G64gat), .B1(new_n722_), .B2(new_n460_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT48), .ZN(new_n729_));
  INV_X1    g528(.A(G64gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n730_), .A3(new_n647_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  INV_X1    g532(.A(new_n722_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n577_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n725_), .A2(new_n733_), .A3(new_n577_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT109), .ZN(G1334gat));
  NOR2_X1   g539(.A1(new_n659_), .A2(G78gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT111), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n725_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G78gat), .B1(new_n722_), .B2(new_n659_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT110), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(KEYINPUT50), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(KEYINPUT50), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(G1335gat));
  INV_X1    g547(.A(new_n363_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n340_), .A2(new_n245_), .A3(new_n749_), .A4(new_n341_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n666_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n602_), .B1(new_n752_), .B2(new_n611_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT112), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n750_), .B(KEYINPUT113), .Z(new_n755_));
  AND3_X1   g554(.A1(new_n681_), .A2(KEYINPUT114), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT114), .B1(new_n681_), .B2(new_n755_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n611_), .A2(new_n602_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n754_), .B1(new_n758_), .B2(new_n759_), .ZN(G1336gat));
  INV_X1    g559(.A(new_n752_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G92gat), .B1(new_n761_), .B2(new_n647_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT115), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n647_), .A2(G92gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n758_), .B2(new_n764_), .ZN(G1337gat));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n257_), .A3(new_n577_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n756_), .A2(new_n757_), .A3(new_n579_), .ZN(new_n767_));
  INV_X1    g566(.A(G99gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n681_), .A2(new_n663_), .A3(new_n755_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G106gat), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT116), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n774_), .A3(G106gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(KEYINPUT52), .A3(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n761_), .A2(new_n258_), .A3(new_n663_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n772_), .A2(KEYINPUT116), .A3(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n776_), .A2(new_n782_), .A3(new_n777_), .A4(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1339gat));
  INV_X1    g583(.A(G113gat), .ZN(new_n785_));
  INV_X1    g584(.A(new_n349_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n351_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n350_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n354_), .A2(new_n349_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n361_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n356_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n361_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n338_), .A2(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n325_), .A2(new_n327_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(KEYINPUT55), .C1(new_n331_), .C2(new_n330_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n332_), .B2(new_n328_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n317_), .B1(new_n328_), .B2(new_n321_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n337_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT56), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n333_), .A2(new_n337_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(new_n804_), .A3(new_n337_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n802_), .A2(new_n803_), .A3(new_n363_), .A4(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n794_), .A2(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n807_), .A2(KEYINPUT57), .A3(new_n640_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT57), .B1(new_n807_), .B2(new_n640_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n673_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n800_), .A2(new_n804_), .A3(new_n337_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n804_), .B1(new_n800_), .B2(new_n337_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n803_), .A4(new_n793_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n802_), .A2(new_n803_), .A3(new_n793_), .A4(new_n805_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT117), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT118), .B1(new_n817_), .B2(new_n819_), .ZN(new_n821_));
  OR3_X1    g620(.A1(new_n817_), .A2(KEYINPUT118), .A3(new_n819_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n811_), .A2(new_n820_), .A3(new_n821_), .A4(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n810_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n810_), .A2(new_n823_), .A3(KEYINPUT119), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n245_), .A3(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n314_), .A2(new_n749_), .A3(new_n342_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT54), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n611_), .A2(new_n647_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n663_), .A2(new_n579_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n785_), .B1(new_n836_), .B2(new_n749_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n824_), .A2(new_n245_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n830_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n835_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n749_), .A2(new_n785_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n834_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n841_), .B(new_n842_), .C1(new_n843_), .C2(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n837_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n837_), .A2(KEYINPUT120), .A3(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1340gat));
  XOR2_X1   g648(.A(KEYINPUT121), .B(G120gat), .Z(new_n850_));
  NAND2_X1  g649(.A1(new_n836_), .A2(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n841_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n852_), .B2(new_n342_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n850_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n342_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n843_), .B(new_n855_), .C1(KEYINPUT60), .C2(new_n854_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1341gat));
  AOI21_X1  g656(.A(G127gat), .B1(new_n843_), .B2(new_n244_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n858_), .A2(KEYINPUT122), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n851_), .A2(G127gat), .A3(new_n244_), .A4(new_n841_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(KEYINPUT122), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(G1342gat));
  AOI21_X1  g661(.A(G134gat), .B1(new_n843_), .B2(new_n641_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n852_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n811_), .A2(G134gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1343gat));
  NOR2_X1   g665(.A1(new_n659_), .A2(new_n577_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n832_), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n868_), .B(new_n869_), .C1(new_n828_), .C2(new_n830_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n363_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g671(.A(new_n342_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT123), .B(G148gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1345gat));
  NAND3_X1  g675(.A1(new_n870_), .A2(new_n491_), .A3(new_n244_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n831_), .A2(new_n867_), .A3(new_n244_), .A4(new_n832_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G155gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n877_), .A2(new_n879_), .A3(new_n881_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1346gat));
  AOI21_X1  g684(.A(G162gat), .B1(new_n870_), .B2(new_n641_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n673_), .A2(new_n492_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n870_), .B2(new_n887_), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n637_), .A2(new_n460_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n830_), .B2(new_n838_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n891_), .A2(new_n363_), .A3(new_n387_), .A4(new_n833_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n833_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n749_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n894_), .B2(new_n384_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT62), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n384_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(KEYINPUT62), .B2(new_n897_), .ZN(G1348gat));
  INV_X1    g697(.A(new_n893_), .ZN(new_n899_));
  AOI21_X1  g698(.A(G176gat), .B1(new_n899_), .B2(new_n873_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n890_), .A2(new_n579_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n663_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n902_), .A2(G176gat), .A3(new_n873_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(G1349gat));
  NOR3_X1   g703(.A1(new_n893_), .A2(new_n406_), .A3(new_n245_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n902_), .A2(new_n244_), .A3(new_n901_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n389_), .B2(new_n906_), .ZN(G1350gat));
  NOR2_X1   g706(.A1(new_n893_), .A2(new_n673_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n641_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n909_));
  OAI22_X1  g708(.A1(new_n908_), .A2(new_n390_), .B1(new_n893_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  OAI221_X1 g711(.A(KEYINPUT125), .B1(new_n893_), .B2(new_n909_), .C1(new_n908_), .C2(new_n390_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1351gat));
  AOI21_X1  g713(.A(new_n868_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n915_), .A2(new_n889_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n363_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n873_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT126), .B(G204gat), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n919_), .B(new_n921_), .ZN(G1353gat));
  NAND2_X1  g721(.A1(new_n916_), .A2(new_n244_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n923_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT63), .B(G211gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n916_), .A2(new_n244_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1354gat));
  NAND3_X1  g726(.A1(new_n915_), .A2(new_n641_), .A3(new_n889_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(G218gat), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n915_), .A2(KEYINPUT127), .A3(new_n641_), .A4(new_n889_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n916_), .A2(G218gat), .A3(new_n811_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1355gat));
endmodule


