//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT71), .B(G1gat), .ZN(new_n206_));
  INV_X1    g005(.A(G8gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT72), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n213_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G29gat), .B(G36gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n219_), .B(KEYINPUT15), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n214_), .A2(new_n215_), .A3(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n219_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n214_), .A2(new_n215_), .A3(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n221_), .B1(new_n220_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n205_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n220_), .A2(new_n227_), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n224_), .B(new_n204_), .C1(new_n230_), .C2(new_n221_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT87), .Z(new_n237_));
  AND2_X1   g036(.A1(G141gat), .A2(G148gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G141gat), .A2(G148gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240_));
  AOI22_X1  g039(.A1(KEYINPUT2), .A2(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(KEYINPUT2), .B2(new_n238_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n234_), .B(new_n235_), .C1(new_n237_), .C2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n238_), .A2(new_n239_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT86), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n245_), .B1(new_n234_), .B2(KEYINPUT1), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n234_), .A2(KEYINPUT1), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n235_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n234_), .A2(new_n245_), .A3(KEYINPUT1), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n244_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n243_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G127gat), .B(G134gat), .Z(new_n252_));
  XOR2_X1   g051(.A(G113gat), .B(G120gat), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n243_), .A2(new_n254_), .A3(new_n250_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(KEYINPUT4), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G225gat), .A2(G233gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n251_), .A2(new_n261_), .A3(new_n255_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n258_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n256_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G1gat), .B(G29gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(G85gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT0), .B(G57gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n263_), .A2(new_n264_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G78gat), .B(G106gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n251_), .A2(KEYINPUT29), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G228gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT89), .B(G197gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G204gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT90), .ZN(new_n279_));
  INV_X1    g078(.A(G204gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(G197gat), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n279_), .A3(G204gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n283_), .A3(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(KEYINPUT91), .B(KEYINPUT21), .Z(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n277_), .A2(new_n280_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n285_), .B1(G197gat), .B2(G204gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n284_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n287_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n275_), .A2(new_n276_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n276_), .B1(new_n275_), .B2(new_n294_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n274_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT92), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT92), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n300_), .B(new_n274_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT28), .B1(new_n251_), .B2(KEYINPUT29), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n251_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G22gat), .B(G50gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n303_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  OR3_X1    g106(.A1(new_n251_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n305_), .B1(new_n308_), .B2(new_n302_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n297_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n274_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n295_), .A3(new_n312_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n299_), .A2(new_n301_), .A3(new_n310_), .A4(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n298_), .A2(new_n313_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT88), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n306_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n308_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT88), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n315_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n273_), .B1(new_n314_), .B2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G8gat), .B(G36gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT18), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G64gat), .B(G92gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT26), .B(G190gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT25), .B(G183gat), .Z(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT23), .ZN(new_n333_));
  OR2_X1    g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT24), .A3(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n334_), .A2(KEYINPUT24), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n331_), .A2(new_n333_), .A3(new_n336_), .A4(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n333_), .B1(G183gat), .B2(G190gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(KEYINPUT22), .B(G169gat), .Z(new_n340_));
  OAI211_X1 g139(.A(new_n339_), .B(new_n335_), .C1(G176gat), .C2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n294_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n345_));
  INV_X1    g144(.A(G183gat), .ZN(new_n346_));
  OR3_X1    g145(.A1(new_n345_), .A2(new_n346_), .A3(KEYINPUT25), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT25), .B1(new_n345_), .B2(new_n346_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n328_), .A3(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n349_), .A2(new_n333_), .A3(new_n336_), .A4(new_n337_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n339_), .A2(new_n335_), .ZN(new_n351_));
  INV_X1    g150(.A(G176gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(G169gat), .B1(KEYINPUT79), .B2(KEYINPUT22), .ZN(new_n353_));
  AND2_X1   g152(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(KEYINPUT77), .A2(G169gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(KEYINPUT77), .A2(G169gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT22), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT78), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(KEYINPUT22), .C1(new_n356_), .C2(new_n357_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n355_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n350_), .B1(new_n351_), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT20), .B1(new_n294_), .B2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n344_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n342_), .A2(new_n294_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT20), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n294_), .B2(new_n363_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n367_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n327_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n368_), .B1(new_n344_), .B2(new_n364_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n370_), .A2(new_n372_), .A3(new_n367_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n326_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(KEYINPUT27), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT95), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT95), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n374_), .A2(new_n380_), .A3(KEYINPUT27), .A4(new_n377_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n326_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n377_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT27), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(KEYINPUT96), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT96), .B1(new_n385_), .B2(new_n386_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n322_), .B(new_n382_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(KEYINPUT32), .B(new_n326_), .C1(new_n369_), .C2(new_n373_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n326_), .A2(KEYINPUT32), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n375_), .A2(new_n376_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n273_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n256_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n395_), .A2(new_n269_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT94), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n258_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n397_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n384_), .B(new_n377_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT33), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n272_), .B(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n394_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n314_), .A2(new_n321_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n390_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n408_));
  INV_X1    g207(.A(G99gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G227gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G71gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n410_), .B(KEYINPUT81), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(G71gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n409_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(G15gat), .B(G43gat), .Z(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(G71gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n412_), .A2(new_n413_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(G99gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n419_), .B1(new_n417_), .B2(new_n422_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n424_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n417_), .A2(new_n422_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n418_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n426_), .B1(new_n430_), .B2(new_n423_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n408_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n427_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n426_), .A3(new_n423_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(KEYINPUT84), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n363_), .A2(KEYINPUT80), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT80), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n350_), .B(new_n437_), .C1(new_n351_), .C2(new_n362_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(KEYINPUT30), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n438_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT30), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n432_), .A2(new_n435_), .A3(new_n439_), .A4(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT84), .B1(new_n433_), .B2(new_n434_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n439_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT31), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n443_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n254_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n443_), .A2(new_n447_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT31), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n255_), .A3(new_n449_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n407_), .A2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n405_), .B(new_n382_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n273_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n452_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n233_), .B1(new_n457_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT13), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(KEYINPUT68), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(KEYINPUT68), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT6), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(G99gat), .A3(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT7), .ZN(new_n473_));
  INV_X1    g272(.A(G106gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n409_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n471_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT65), .B1(new_n476_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  OR2_X1    g280(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT64), .ZN(new_n483_));
  NAND2_X1  g282(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n474_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n477_), .A2(KEYINPUT9), .A3(new_n478_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n478_), .A2(KEYINPUT9), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n488_), .A2(new_n471_), .A3(new_n489_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n480_), .A2(new_n481_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n468_), .A2(new_n470_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n475_), .A2(new_n472_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n479_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT65), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n476_), .A2(KEYINPUT65), .A3(new_n479_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(KEYINPUT8), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n501_));
  XOR2_X1   g300(.A(G71gat), .B(G78gat), .Z(new_n502_));
  OR2_X1    g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n502_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT66), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n499_), .A2(new_n507_), .B1(new_n508_), .B2(KEYINPUT12), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n476_), .A2(KEYINPUT65), .A3(new_n479_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n510_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n487_), .A2(new_n490_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n496_), .B2(KEYINPUT8), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n507_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n491_), .A2(new_n498_), .A3(new_n506_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT66), .B(KEYINPUT12), .Z(new_n517_));
  AOI21_X1  g316(.A(new_n509_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G230gat), .A2(G233gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G120gat), .B(G148gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT5), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G176gat), .B(G204gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT67), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n520_), .A2(new_n522_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n465_), .B(new_n466_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n530_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(KEYINPUT13), .A4(new_n528_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G134gat), .B(G162gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(G190gat), .B(G218gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n539_), .A2(new_n540_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n511_), .A2(new_n513_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n543_), .A2(new_n219_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n544_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n499_), .B2(new_n222_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT70), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n548_), .A2(KEYINPUT70), .A3(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n549_), .ZN(new_n556_));
  OAI22_X1  g355(.A1(new_n499_), .A2(new_n226_), .B1(KEYINPUT35), .B2(new_n546_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n499_), .A2(new_n222_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n557_), .B1(KEYINPUT69), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(KEYINPUT69), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n556_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n541_), .B(new_n542_), .C1(new_n555_), .C2(new_n562_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n548_), .A2(KEYINPUT70), .A3(new_n550_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT70), .B1(new_n548_), .B2(new_n550_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n558_), .A2(KEYINPUT69), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n548_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n549_), .B1(new_n568_), .B2(new_n560_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n566_), .A2(new_n569_), .A3(new_n540_), .A4(new_n539_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n563_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT37), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(G231gat), .ZN(new_n575_));
  INV_X1    g374(.A(G233gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n506_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n575_), .A2(new_n576_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n503_), .B(new_n578_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT73), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT73), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(new_n579_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n216_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n581_), .A2(new_n214_), .A3(new_n215_), .A4(new_n583_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT16), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT74), .B1(new_n587_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n591_), .B(KEYINPUT17), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n585_), .A2(new_n586_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT75), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT75), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n585_), .A2(new_n598_), .A3(new_n586_), .A4(new_n595_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n594_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n594_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT37), .B1(new_n563_), .B2(new_n570_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n536_), .A2(new_n574_), .A3(new_n602_), .A4(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n462_), .A2(KEYINPUT97), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n390_), .A2(new_n406_), .B1(new_n455_), .B2(new_n452_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n458_), .A2(new_n460_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n232_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n608_), .B1(new_n611_), .B2(new_n605_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n607_), .A2(new_n612_), .A3(KEYINPUT98), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n615_), .A2(new_n273_), .A3(new_n206_), .A4(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n600_), .A2(new_n601_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n620_), .A2(new_n535_), .A3(new_n233_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n621_), .B(new_n571_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n459_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n617_), .A2(new_n618_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n619_), .A2(new_n623_), .A3(new_n624_), .ZN(G1324gat));
  XNOR2_X1  g424(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628_));
  INV_X1    g427(.A(new_n377_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n386_), .B1(new_n629_), .B2(new_n383_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n632_), .A2(new_n387_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n633_), .A2(new_n322_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n456_), .ZN(new_n635_));
  OAI22_X1  g434(.A1(new_n634_), .A2(new_n635_), .B1(new_n460_), .B2(new_n458_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n633_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n571_), .A4(new_n621_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(G8gat), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n639_), .B1(new_n638_), .B2(G8gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n628_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n642_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(KEYINPUT100), .A3(new_n640_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n643_), .A2(new_n645_), .A3(KEYINPUT39), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n615_), .A2(new_n207_), .A3(new_n637_), .A4(new_n616_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n628_), .B(new_n648_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n627_), .B1(new_n646_), .B2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n643_), .A2(new_n645_), .A3(KEYINPUT39), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n652_), .A2(new_n649_), .A3(new_n647_), .A4(new_n626_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n622_), .B2(new_n456_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT41), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n613_), .A2(G15gat), .A3(new_n456_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1326gat));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  INV_X1    g458(.A(new_n622_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n405_), .B(KEYINPUT102), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n659_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT42), .Z(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n659_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT103), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n613_), .B2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n571_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n620_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n535_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n462_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G29gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n273_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n674_));
  NOR4_X1   g473(.A1(new_n602_), .A2(new_n535_), .A3(new_n233_), .A4(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n574_), .A2(new_n604_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n676_), .B(new_n677_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n676_), .B1(new_n636_), .B2(new_n677_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT105), .B1(KEYINPUT104), .B2(KEYINPUT44), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n675_), .B(new_n682_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n459_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n673_), .B1(new_n686_), .B2(new_n672_), .ZN(G1328gat));
  INV_X1    g486(.A(G36gat), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n637_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n670_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT45), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n633_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n688_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(KEYINPUT106), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697_));
  OAI221_X1 g496(.A(new_n692_), .B1(new_n697_), .B2(KEYINPUT46), .C1(new_n693_), .C2(new_n688_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1329gat));
  NAND2_X1  g498(.A1(new_n684_), .A2(new_n685_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(G43gat), .A3(new_n635_), .ZN(new_n701_));
  INV_X1    g500(.A(G43gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n670_), .B2(new_n456_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT107), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n701_), .A2(new_n704_), .A3(new_n706_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1330gat));
  AOI21_X1  g509(.A(G50gat), .B1(new_n671_), .B2(new_n661_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n405_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n700_), .B2(new_n713_), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n609_), .A2(new_n610_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(new_n232_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n620_), .A2(new_n573_), .A3(new_n603_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(new_n535_), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(G57gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n273_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n715_), .A2(new_n667_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n536_), .A2(new_n620_), .A3(new_n232_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G57gat), .B1(new_n723_), .B2(new_n459_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n720_), .A2(new_n724_), .ZN(G1332gat));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n718_), .A2(new_n726_), .A3(new_n637_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n721_), .A2(new_n637_), .A3(new_n722_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(G64gat), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n728_), .B2(G64gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT109), .Z(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n723_), .B2(new_n456_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT49), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n635_), .A2(new_n413_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT110), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n718_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1334gat));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  INV_X1    g540(.A(new_n723_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(new_n661_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT50), .Z(new_n744_));
  NAND2_X1  g543(.A1(new_n661_), .A2(new_n741_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT111), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n718_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n747_), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n668_), .A2(new_n536_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n716_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(G85gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n273_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n620_), .A2(new_n535_), .A3(new_n233_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n677_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT43), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n756_), .B2(new_n678_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(new_n273_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n753_), .B1(new_n758_), .B2(new_n752_), .ZN(G1336gat));
  AOI21_X1  g558(.A(G92gat), .B1(new_n751_), .B2(new_n637_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n761_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n637_), .A2(G92gat), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n762_), .A2(new_n763_), .B1(new_n757_), .B2(new_n764_), .ZN(G1337gat));
  NOR2_X1   g564(.A1(new_n485_), .A2(new_n486_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n456_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT113), .B1(new_n751_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  INV_X1    g568(.A(new_n767_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n750_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n757_), .A2(new_n635_), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n768_), .A2(new_n771_), .B1(new_n772_), .B2(new_n409_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n751_), .A2(new_n474_), .A3(new_n712_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n757_), .A2(new_n712_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(G106gat), .ZN(new_n778_));
  AOI211_X1 g577(.A(KEYINPUT52), .B(new_n474_), .C1(new_n757_), .C2(new_n712_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n782_), .B(new_n775_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1339gat));
  NOR3_X1   g583(.A1(new_n637_), .A2(new_n456_), .A3(new_n459_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n520_), .A2(new_n522_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n526_), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n229_), .A2(new_n231_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n518_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n519_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n491_), .A2(new_n498_), .A3(new_n506_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n506_), .B1(new_n491_), .B2(new_n498_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n517_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n508_), .A2(KEYINPUT12), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n514_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n792_), .A2(KEYINPUT55), .A3(new_n519_), .A4(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n792_), .A2(new_n794_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n521_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n521_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n789_), .B(new_n797_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n526_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n526_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n788_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n221_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n220_), .A2(new_n806_), .A3(new_n223_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n205_), .B(new_n807_), .C1(new_n230_), .C2(new_n806_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n231_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n532_), .A2(new_n528_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT116), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n805_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n571_), .A2(KEYINPUT116), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT57), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n816_), .B(new_n813_), .C1(new_n805_), .C2(new_n811_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n786_), .A2(new_n787_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n819_), .A2(new_n231_), .A3(new_n808_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(KEYINPUT58), .C1(new_n804_), .C2(new_n803_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n820_), .B1(new_n804_), .B2(new_n803_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n802_), .A2(new_n526_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n526_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n831_), .A2(KEYINPUT117), .A3(KEYINPUT58), .A4(new_n820_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n823_), .A2(new_n677_), .A3(new_n826_), .A4(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n602_), .B1(new_n818_), .B2(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n605_), .B2(new_n232_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(KEYINPUT114), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n717_), .A2(new_n233_), .A3(new_n536_), .A4(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n405_), .B(new_n785_), .C1(new_n834_), .C2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n232_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n812_), .A2(new_n814_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n816_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n812_), .A2(KEYINPUT57), .A3(new_n814_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n833_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n840_), .B1(new_n848_), .B2(new_n620_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n712_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(KEYINPUT118), .A3(KEYINPUT59), .A4(new_n785_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n841_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n233_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n844_), .B1(new_n855_), .B2(new_n843_), .ZN(G1340gat));
  XNOR2_X1  g655(.A(KEYINPUT119), .B(G120gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT60), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n535_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT120), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n842_), .B(new_n861_), .C1(new_n860_), .C2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n536_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n857_), .ZN(G1341gat));
  INV_X1    g665(.A(G127gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n842_), .A2(new_n867_), .A3(new_n602_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n620_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1342gat));
  AOI21_X1  g669(.A(G134gat), .B1(new_n842_), .B2(new_n667_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n851_), .A2(new_n854_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT121), .B(G134gat), .Z(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n574_), .B2(new_n604_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n871_), .B1(new_n872_), .B2(new_n874_), .ZN(G1343gat));
  NOR4_X1   g674(.A1(new_n635_), .A2(new_n637_), .A3(new_n405_), .A4(new_n459_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n849_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n232_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n535_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g681(.A1(new_n848_), .A2(new_n620_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n840_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n602_), .A3(new_n876_), .ZN(new_n886_));
  XOR2_X1   g685(.A(KEYINPUT61), .B(G155gat), .Z(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n889_));
  INV_X1    g688(.A(new_n887_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n878_), .A2(new_n602_), .A3(new_n890_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n888_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n889_), .B1(new_n888_), .B2(new_n891_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1346gat));
  INV_X1    g693(.A(G162gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n878_), .A2(new_n895_), .A3(new_n667_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n878_), .A2(new_n677_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n895_), .ZN(G1347gat));
  OR2_X1    g697(.A1(new_n460_), .A2(new_n633_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n661_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n232_), .B(new_n900_), .C1(new_n834_), .C2(new_n840_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n902_));
  INV_X1    g701(.A(new_n340_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n885_), .A2(new_n903_), .A3(new_n232_), .A4(new_n900_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(KEYINPUT62), .B1(new_n901_), .B2(G169gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT124), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n901_), .A2(G169gat), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n910_), .A2(new_n911_), .A3(new_n904_), .A4(new_n902_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n907_), .A2(new_n912_), .ZN(G1348gat));
  NAND2_X1  g712(.A1(new_n885_), .A2(new_n900_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(G176gat), .B1(new_n915_), .B2(new_n535_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n849_), .A2(new_n712_), .A3(new_n899_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n536_), .A2(new_n352_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(G1349gat));
  NOR4_X1   g718(.A1(new_n849_), .A2(new_n712_), .A3(new_n620_), .A4(new_n899_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n602_), .A2(new_n330_), .ZN(new_n921_));
  OAI22_X1  g720(.A1(new_n920_), .A2(G183gat), .B1(new_n914_), .B2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT125), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924_));
  OAI221_X1 g723(.A(new_n924_), .B1(new_n914_), .B2(new_n921_), .C1(new_n920_), .C2(G183gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n915_), .A2(new_n328_), .A3(new_n667_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n914_), .B1(new_n574_), .B2(new_n604_), .ZN(new_n928_));
  INV_X1    g727(.A(G190gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(G1351gat));
  AND3_X1   g729(.A1(new_n637_), .A2(new_n456_), .A3(new_n322_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n885_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n232_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n535_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G204gat), .ZN(G1353gat));
  AND3_X1   g735(.A1(new_n885_), .A2(new_n602_), .A3(new_n931_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT63), .B(G211gat), .Z(new_n938_));
  AOI21_X1  g737(.A(KEYINPUT126), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n885_), .A2(new_n602_), .A3(new_n931_), .A4(new_n938_), .ZN(new_n940_));
  OR2_X1    g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n937_), .B2(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n939_), .B1(KEYINPUT126), .B2(new_n942_), .ZN(G1354gat));
  NAND2_X1  g742(.A1(new_n932_), .A2(new_n667_), .ZN(new_n944_));
  XOR2_X1   g743(.A(KEYINPUT127), .B(G218gat), .Z(new_n945_));
  AOI21_X1  g744(.A(new_n945_), .B1(new_n574_), .B2(new_n604_), .ZN(new_n946_));
  AOI22_X1  g745(.A1(new_n944_), .A2(new_n945_), .B1(new_n932_), .B2(new_n946_), .ZN(G1355gat));
endmodule


