//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n839_, new_n841_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT6), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT66), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n208_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n210_), .B(new_n211_), .C1(new_n206_), .C2(KEYINPUT66), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n205_), .A2(new_n207_), .A3(new_n209_), .A4(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT67), .B(KEYINPUT8), .Z(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT67), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .A4(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n215_), .A2(KEYINPUT65), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT9), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(KEYINPUT9), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n214_), .A3(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n204_), .B(KEYINPUT6), .Z(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT10), .B(G99gat), .Z(new_n228_));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n211_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT10), .B(G99gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT64), .B1(new_n231_), .B2(G106gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n227_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n218_), .A2(new_n222_), .B1(new_n226_), .B2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G57gat), .B(G64gat), .Z(new_n235_));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238_));
  XOR2_X1   g037(.A(G71gat), .B(G78gat), .Z(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n238_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n242_));
  OAI22_X1  g041(.A1(new_n241_), .A2(new_n242_), .B1(new_n236_), .B2(new_n235_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n235_), .A2(new_n236_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n240_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n234_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT69), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n234_), .A2(new_n247_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n234_), .A2(new_n247_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n203_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n218_), .A2(new_n222_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n233_), .A2(new_n226_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT70), .B1(new_n233_), .B2(new_n226_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n256_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n261_), .A2(KEYINPUT12), .A3(new_n246_), .A4(new_n243_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(new_n234_), .B2(new_n247_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n262_), .A2(new_n202_), .A3(new_n248_), .A4(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n255_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT5), .B(G176gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G204gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(G120gat), .B(G148gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(KEYINPUT71), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT13), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT13), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G15gat), .B(G22gat), .ZN(new_n278_));
  INV_X1    g077(.A(G1gat), .ZN(new_n279_));
  INV_X1    g078(.A(G8gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT14), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G1gat), .B(G8gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G29gat), .B(G36gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G43gat), .B(G50gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT78), .Z(new_n290_));
  NAND2_X1  g089(.A1(G229gat), .A2(G233gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n287_), .B(KEYINPUT15), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n284_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n290_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n284_), .A2(new_n288_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT79), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n290_), .A2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n295_), .B1(new_n298_), .B2(new_n291_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G113gat), .B(G141gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G169gat), .B(G197gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n301_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n277_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G22gat), .B(G50gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(G211gat), .B(G218gat), .Z(new_n309_));
  XOR2_X1   g108(.A(G197gat), .B(G204gat), .Z(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT21), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT88), .ZN(new_n312_));
  OR3_X1    g111(.A1(new_n310_), .A2(KEYINPUT87), .A3(KEYINPUT21), .ZN(new_n313_));
  INV_X1    g112(.A(new_n309_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT21), .B1(new_n310_), .B2(KEYINPUT87), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n318_));
  OR4_X1    g117(.A1(new_n318_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  INV_X1    g119(.A(G141gat), .ZN(new_n321_));
  INV_X1    g120(.A(G148gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n320_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  OAI22_X1  g122(.A1(new_n318_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n319_), .A2(new_n323_), .A3(new_n324_), .A4(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  INV_X1    g126(.A(G155gat), .ZN(new_n328_));
  INV_X1    g127(.A(G162gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(KEYINPUT83), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT83), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(G155gat), .B2(G162gat), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n326_), .A2(new_n327_), .A3(new_n330_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(KEYINPUT1), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(new_n334_), .A3(new_n332_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT84), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n327_), .A2(KEYINPUT1), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT84), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n330_), .A2(new_n334_), .A3(new_n332_), .A4(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n341_));
  XOR2_X1   g140(.A(G141gat), .B(G148gat), .Z(new_n342_));
  AND3_X1   g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n333_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n317_), .B1(new_n345_), .B2(KEYINPUT29), .ZN(new_n346_));
  INV_X1    g145(.A(G228gat), .ZN(new_n347_));
  INV_X1    g146(.A(G233gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  AOI211_X1 g150(.A(new_n349_), .B(new_n317_), .C1(KEYINPUT29), .C2(new_n345_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n308_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n345_), .A2(KEYINPUT29), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G78gat), .B(G106gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT28), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n354_), .B(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n345_), .A2(KEYINPUT29), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n312_), .A2(new_n316_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n349_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n346_), .A2(new_n350_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n308_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n353_), .A2(new_n358_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n358_), .B1(new_n365_), .B2(new_n353_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(G71gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(G183gat), .A3(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n375_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT81), .B1(new_n375_), .B2(KEYINPUT23), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n374_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT25), .B(G183gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT26), .B(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G169gat), .ZN(new_n382_));
  INV_X1    g181(.A(G176gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n384_), .A2(KEYINPUT24), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(KEYINPUT24), .A3(new_n386_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n378_), .A2(new_n381_), .A3(new_n385_), .A4(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n386_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT22), .B(G169gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n390_), .B2(new_n383_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n375_), .A2(KEYINPUT23), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n392_), .A2(new_n374_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n391_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT30), .B(G99gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n388_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n388_), .B2(new_n395_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n372_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n388_), .A2(new_n395_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n396_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n372_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(new_n397_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G15gat), .B(G43gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n400_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n406_), .B1(new_n400_), .B2(new_n405_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n369_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n400_), .A2(new_n405_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n406_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(KEYINPUT82), .A3(new_n407_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G127gat), .B(G134gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G113gat), .B(G120gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT31), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n410_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n418_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n369_), .B(new_n420_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n368_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n417_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n345_), .A2(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n417_), .B(new_n333_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(KEYINPUT4), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT91), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n425_), .A2(KEYINPUT4), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n425_), .A2(KEYINPUT91), .A3(KEYINPUT4), .A4(new_n426_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n429_), .A2(new_n431_), .A3(new_n432_), .A4(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n425_), .A2(new_n426_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n430_), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT92), .B(KEYINPUT0), .Z(new_n437_));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G57gat), .B(G85gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n434_), .A2(new_n436_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT94), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n443_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n434_), .A2(KEYINPUT33), .A3(new_n436_), .A4(new_n441_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n441_), .B1(new_n435_), .B2(new_n431_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n429_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(new_n449_), .B2(new_n431_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n381_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n451_), .A2(new_n393_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n378_), .B1(G183gat), .B2(G190gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n391_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n360_), .A2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n456_), .B(KEYINPUT20), .C1(new_n401_), .C2(new_n360_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G226gat), .A2(G233gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n458_), .B(KEYINPUT19), .Z(new_n459_));
  XOR2_X1   g258(.A(new_n459_), .B(KEYINPUT89), .Z(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT90), .B(KEYINPUT18), .Z(new_n462_));
  XNOR2_X1  g261(.A(G8gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G64gat), .B(G92gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n360_), .A2(new_n401_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n312_), .A2(new_n316_), .A3(new_n454_), .A4(new_n452_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n468_), .A2(KEYINPUT20), .A3(new_n459_), .A4(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n461_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n467_), .B1(new_n461_), .B2(new_n470_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n447_), .A2(new_n450_), .A3(new_n473_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n445_), .A2(new_n446_), .A3(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n468_), .A2(KEYINPUT20), .A3(new_n469_), .ZN(new_n476_));
  OAI22_X1  g275(.A1(new_n476_), .A2(new_n459_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n467_), .A2(KEYINPUT32), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n459_), .A2(new_n476_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT32), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n480_), .B1(new_n481_), .B2(new_n466_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n442_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n441_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n479_), .B(new_n482_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n423_), .B1(new_n475_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n422_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n358_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n365_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n364_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n419_), .A2(new_n421_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n353_), .A2(new_n358_), .A3(new_n365_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n488_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT27), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT96), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT96), .B(new_n497_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT95), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(new_n480_), .B2(new_n467_), .ZN(new_n503_));
  AND4_X1   g302(.A1(new_n502_), .A2(new_n461_), .A3(new_n467_), .A4(new_n470_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n497_), .B1(new_n477_), .B2(new_n466_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n500_), .A2(new_n501_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n483_), .A2(new_n484_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n496_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n307_), .B1(new_n487_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n257_), .B(new_n258_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n292_), .B1(new_n514_), .B2(new_n256_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n234_), .A2(new_n287_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT35), .B(new_n513_), .C1(new_n515_), .C2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n261_), .A2(new_n293_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n513_), .A2(KEYINPUT35), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n513_), .A2(KEYINPUT35), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .A4(new_n516_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT74), .ZN(new_n524_));
  XOR2_X1   g323(.A(G190gat), .B(G218gat), .Z(new_n525_));
  XNOR2_X1  g324(.A(G134gat), .B(G162gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT36), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT74), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n518_), .A2(new_n529_), .A3(new_n522_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT75), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n523_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT75), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n524_), .A2(new_n537_), .A3(new_n528_), .A4(new_n530_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT76), .B(KEYINPUT37), .Z(new_n539_));
  NAND4_X1  g338(.A1(new_n532_), .A2(new_n536_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n528_), .A2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n528_), .A2(new_n541_), .ZN(new_n543_));
  AOI211_X1 g342(.A(new_n542_), .B(new_n543_), .C1(new_n518_), .C2(new_n522_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT37), .B1(new_n544_), .B2(new_n535_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n284_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n247_), .ZN(new_n549_));
  XOR2_X1   g348(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n550_));
  XNOR2_X1  g349(.A(G127gat), .B(G155gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G183gat), .B(G211gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT17), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n554_), .B(KEYINPUT17), .Z(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n549_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n546_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n510_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n508_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n279_), .A3(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT97), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT38), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n532_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT98), .Z(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n487_), .B2(new_n509_), .ZN(new_n569_));
  AND4_X1   g368(.A1(new_n558_), .A2(new_n569_), .A3(new_n306_), .A4(new_n277_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n279_), .B1(new_n570_), .B2(new_n563_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT99), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(G1324gat));
  INV_X1    g372(.A(new_n507_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n280_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT39), .Z(new_n576_));
  NAND3_X1  g375(.A1(new_n562_), .A2(new_n280_), .A3(new_n574_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g378(.A(G15gat), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n570_), .B2(new_n422_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT41), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n562_), .A2(new_n580_), .A3(new_n422_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(G1326gat));
  INV_X1    g383(.A(G22gat), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n570_), .B2(new_n368_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT42), .Z(new_n587_));
  NAND3_X1  g386(.A1(new_n562_), .A2(new_n585_), .A3(new_n368_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(G1327gat));
  INV_X1    g388(.A(KEYINPUT43), .ZN(new_n590_));
  INV_X1    g389(.A(new_n368_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n493_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n474_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n442_), .A2(new_n444_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT94), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n592_), .B1(new_n597_), .B2(new_n485_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n496_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n590_), .B(new_n546_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n487_), .A2(new_n509_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n603_), .A2(KEYINPUT100), .A3(new_n590_), .A4(new_n546_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n546_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT43), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n307_), .A2(new_n558_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT44), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n607_), .A2(KEYINPUT44), .A3(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G29gat), .B1(new_n613_), .B2(new_n508_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n568_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(new_n558_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n510_), .A2(new_n616_), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n617_), .A2(G29gat), .A3(new_n508_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(G1328gat));
  NAND3_X1  g418(.A1(new_n611_), .A2(new_n574_), .A3(new_n612_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n611_), .A2(KEYINPUT101), .A3(new_n574_), .A4(new_n612_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(G36gat), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT102), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n622_), .A2(new_n626_), .A3(G36gat), .A4(new_n623_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n617_), .A2(G36gat), .A3(new_n507_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT46), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(KEYINPUT46), .A3(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1329gat));
  OAI21_X1  g435(.A(G43gat), .B1(new_n613_), .B2(new_n493_), .ZN(new_n637_));
  OR3_X1    g436(.A1(new_n617_), .A2(G43gat), .A3(new_n493_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(G1330gat));
  OAI21_X1  g440(.A(G50gat), .B1(new_n613_), .B2(new_n591_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n617_), .A2(G50gat), .A3(new_n591_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1331gat));
  NOR2_X1   g443(.A1(new_n277_), .A2(new_n306_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(new_n603_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n560_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT105), .Z(new_n648_));
  AOI21_X1  g447(.A(G57gat), .B1(new_n648_), .B2(new_n563_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n569_), .A2(new_n558_), .A3(new_n645_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(new_n563_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n649_), .B1(G57gat), .B2(new_n651_), .ZN(G1332gat));
  INV_X1    g451(.A(G64gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n650_), .B2(new_n574_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT48), .Z(new_n655_));
  NAND3_X1  g454(.A1(new_n648_), .A2(new_n653_), .A3(new_n574_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1333gat));
  AOI21_X1  g456(.A(new_n371_), .B1(new_n650_), .B2(new_n422_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT49), .Z(new_n659_));
  NAND3_X1  g458(.A1(new_n648_), .A2(new_n371_), .A3(new_n422_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1334gat));
  INV_X1    g460(.A(G78gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n650_), .B2(new_n368_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT50), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n648_), .A2(new_n662_), .A3(new_n368_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1335gat));
  INV_X1    g465(.A(G85gat), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n646_), .A2(new_n616_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(new_n508_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT106), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n607_), .A2(new_n559_), .A3(new_n645_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n508_), .A2(new_n667_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT107), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(new_n671_), .B2(new_n673_), .ZN(G1336gat));
  NOR3_X1   g473(.A1(new_n668_), .A2(G92gat), .A3(new_n507_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n671_), .A2(new_n574_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(G92gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT108), .ZN(G1337gat));
  NOR3_X1   g477(.A1(new_n668_), .A2(new_n231_), .A3(new_n493_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n671_), .A2(new_n422_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(G99gat), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g481(.A(KEYINPUT52), .ZN(new_n683_));
  INV_X1    g482(.A(new_n671_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G106gat), .B1(new_n684_), .B2(new_n591_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(KEYINPUT109), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(KEYINPUT109), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n685_), .A2(KEYINPUT109), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n685_), .A2(KEYINPUT109), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(KEYINPUT52), .A3(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n646_), .A2(new_n616_), .A3(new_n211_), .A4(new_n368_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n688_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT53), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT53), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n688_), .A2(new_n691_), .A3(new_n695_), .A4(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1339gat));
  INV_X1    g496(.A(KEYINPUT57), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n291_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n700_));
  MUX2_X1   g499(.A(new_n299_), .B(new_n700_), .S(new_n304_), .Z(new_n701_));
  NAND2_X1  g500(.A1(new_n274_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT115), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT115), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n274_), .A2(new_n701_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT55), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n265_), .A2(KEYINPUT111), .A3(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT111), .B1(new_n265_), .B2(new_n707_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n262_), .A2(new_n264_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n253_), .B2(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n252_), .A2(KEYINPUT112), .A3(new_n264_), .A4(new_n262_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n203_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(new_n265_), .B2(new_n707_), .ZN(new_n717_));
  OR3_X1    g516(.A1(new_n265_), .A2(new_n716_), .A3(new_n707_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n710_), .A2(new_n715_), .A3(new_n717_), .A4(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT56), .B1(new_n719_), .B2(new_n272_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(KEYINPUT114), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(KEYINPUT56), .A3(new_n272_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n305_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n271_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n720_), .B2(KEYINPUT114), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n706_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n698_), .B1(new_n726_), .B2(new_n568_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT116), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n720_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n722_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n725_), .A3(new_n306_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n703_), .A3(new_n705_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(KEYINPUT57), .A3(new_n615_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT117), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n730_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n720_), .A2(KEYINPUT117), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n722_), .A3(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n739_), .A2(KEYINPUT58), .A3(new_n271_), .A4(new_n701_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT58), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n720_), .A2(KEYINPUT117), .ZN(new_n742_));
  AOI211_X1 g541(.A(new_n736_), .B(KEYINPUT56), .C1(new_n719_), .C2(new_n272_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n722_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n271_), .A2(new_n701_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n741_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n740_), .A2(new_n747_), .A3(new_n546_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT116), .B(new_n698_), .C1(new_n726_), .C2(new_n568_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n729_), .A2(new_n735_), .A3(new_n748_), .A4(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n559_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n560_), .A2(new_n305_), .A3(new_n277_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n752_), .B(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n751_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n574_), .A2(new_n508_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(new_n488_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G113gat), .B1(new_n762_), .B2(new_n306_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(KEYINPUT59), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n748_), .A2(new_n735_), .A3(new_n727_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n755_), .B1(new_n765_), .B2(new_n559_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n760_), .A3(new_n768_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n764_), .A2(G113gat), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n763_), .B1(new_n770_), .B2(new_n306_), .ZN(G1340gat));
  NAND2_X1  g570(.A1(new_n764_), .A2(new_n769_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G120gat), .B1(new_n772_), .B2(new_n277_), .ZN(new_n773_));
  INV_X1    g572(.A(G120gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n277_), .B2(KEYINPUT60), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n774_), .A2(KEYINPUT60), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n757_), .A2(new_n760_), .A3(new_n775_), .A4(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT119), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n773_), .A2(new_n778_), .ZN(G1341gat));
  AOI21_X1  g578(.A(G127gat), .B1(new_n762_), .B2(new_n558_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n764_), .A2(G127gat), .A3(new_n769_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n558_), .ZN(G1342gat));
  INV_X1    g581(.A(G134gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n761_), .B2(new_n615_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n764_), .A2(G134gat), .A3(new_n546_), .A4(new_n769_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT120), .B(new_n783_), .C1(new_n761_), .C2(new_n615_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(G1343gat));
  AOI21_X1  g588(.A(new_n755_), .B1(new_n750_), .B2(new_n559_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(new_n495_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n306_), .A3(new_n758_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT121), .B(G141gat), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1344gat));
  OR2_X1    g593(.A1(new_n790_), .A2(new_n495_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n795_), .A2(new_n277_), .A3(new_n759_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(new_n322_), .ZN(G1345gat));
  NAND3_X1  g596(.A1(new_n791_), .A2(new_n558_), .A3(new_n758_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(KEYINPUT61), .B(G155gat), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(G1346gat));
  NOR2_X1   g599(.A1(new_n795_), .A2(new_n759_), .ZN(new_n801_));
  AOI21_X1  g600(.A(G162gat), .B1(new_n801_), .B2(new_n568_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n546_), .A2(G162gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(new_n803_), .ZN(G1347gat));
  XOR2_X1   g603(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(KEYINPUT123), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(KEYINPUT123), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n507_), .A2(new_n563_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(new_n493_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR4_X1   g612(.A1(new_n766_), .A2(new_n368_), .A3(new_n305_), .A4(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n808_), .B(new_n809_), .C1(new_n814_), .C2(new_n382_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n390_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n767_), .A2(new_n591_), .A3(new_n306_), .A4(new_n812_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(G169gat), .A3(new_n807_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n815_), .A2(new_n816_), .A3(KEYINPUT124), .A4(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1348gat));
  NOR3_X1   g622(.A1(new_n766_), .A2(new_n368_), .A3(new_n813_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n277_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G176gat), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n790_), .A2(new_n368_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n813_), .A2(new_n383_), .A3(new_n277_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(G1349gat));
  INV_X1    g628(.A(new_n379_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n824_), .A2(new_n558_), .A3(new_n830_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n831_), .A2(KEYINPUT125), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(KEYINPUT125), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n813_), .A2(new_n559_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G183gat), .B1(new_n827_), .B2(new_n834_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n832_), .A2(new_n833_), .A3(new_n835_), .ZN(G1350gat));
  NAND3_X1  g635(.A1(new_n824_), .A2(new_n568_), .A3(new_n380_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n824_), .A2(new_n546_), .ZN(new_n838_));
  INV_X1    g637(.A(G190gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(G1351gat));
  NAND3_X1  g639(.A1(new_n791_), .A2(new_n306_), .A3(new_n810_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g641(.A1(new_n791_), .A2(new_n825_), .A3(new_n810_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G204gat), .ZN(G1353gat));
  NOR4_X1   g643(.A1(new_n790_), .A2(new_n559_), .A3(new_n495_), .A4(new_n811_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT63), .ZN(new_n846_));
  INV_X1    g645(.A(G211gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n847_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n845_), .A2(new_n848_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT126), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT126), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n845_), .A2(new_n853_), .A3(new_n848_), .A4(new_n850_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n845_), .A2(new_n848_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n852_), .A2(new_n854_), .A3(new_n855_), .ZN(G1354gat));
  NOR2_X1   g655(.A1(new_n795_), .A2(new_n811_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G218gat), .B1(new_n857_), .B2(new_n568_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n546_), .A2(G218gat), .ZN(new_n859_));
  XOR2_X1   g658(.A(new_n859_), .B(KEYINPUT127), .Z(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n857_), .B2(new_n860_), .ZN(G1355gat));
endmodule


