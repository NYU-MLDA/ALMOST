//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n204_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT83), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G190gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT23), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT83), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n204_), .A2(new_n218_), .A3(new_n208_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n210_), .A2(new_n216_), .A3(new_n217_), .A4(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n207_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT22), .B(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n215_), .A2(KEYINPUT84), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT84), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n216_), .B2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n224_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n220_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231_));
  INV_X1    g030(.A(G204gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(G197gat), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n231_), .B(KEYINPUT21), .C1(KEYINPUT93), .C2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G197gat), .B(G204gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n234_), .A2(new_n235_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n231_), .A2(KEYINPUT21), .ZN(new_n238_));
  NOR3_X1   g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT20), .B1(new_n230_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT97), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n227_), .B1(KEYINPUT98), .B2(new_n209_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n243_), .B(new_n217_), .C1(KEYINPUT98), .C2(new_n209_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n216_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n224_), .B1(new_n245_), .B2(new_n228_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n239_), .ZN(new_n248_));
  OAI211_X1 g047(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n230_), .C2(new_n239_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n242_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G226gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT19), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT96), .Z(new_n253_));
  NAND2_X1  g052(.A1(new_n230_), .A2(new_n239_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n254_), .B(KEYINPUT20), .C1(new_n247_), .C2(new_n239_), .ZN(new_n255_));
  OAI22_X1  g054(.A1(new_n250_), .A2(new_n253_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT18), .B(G64gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G92gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n256_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT27), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n242_), .A2(new_n253_), .A3(new_n248_), .A4(new_n249_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n255_), .A2(new_n252_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n260_), .B(KEYINPUT101), .Z(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n268_), .B(KEYINPUT27), .C1(new_n256_), .C2(new_n260_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT87), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(G43gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT30), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n230_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G43gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G15gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G71gat), .B(G99gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  AND3_X1   g080(.A1(new_n273_), .A2(new_n277_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n273_), .B2(new_n277_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n271_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n273_), .A2(new_n277_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n281_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n273_), .A2(new_n277_), .A3(new_n281_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(KEYINPUT87), .A3(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT85), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT86), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G113gat), .B(G120gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n292_), .B(new_n294_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(new_n293_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT31), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n284_), .A2(new_n289_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n298_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n271_), .B(new_n300_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT88), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT1), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n305_), .A2(KEYINPUT1), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G141gat), .ZN(new_n309_));
  INV_X1    g108(.A(G148gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n316_), .A2(new_n318_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n304_), .B(new_n305_), .C1(new_n321_), .C2(KEYINPUT89), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(KEYINPUT89), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(KEYINPUT90), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT90), .ZN(new_n326_));
  INV_X1    g125(.A(new_n324_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(new_n322_), .B2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n314_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n239_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT92), .ZN(new_n332_));
  INV_X1    g131(.A(G228gat), .ZN(new_n333_));
  INV_X1    g132(.A(G233gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT92), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n336_), .B(new_n239_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n332_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n335_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G78gat), .B(G106gat), .Z(new_n340_));
  NOR3_X1   g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT95), .ZN(new_n342_));
  INV_X1    g141(.A(new_n339_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n340_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n332_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT95), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n329_), .A2(new_n330_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n349_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G22gat), .B(G50gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n340_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n342_), .A2(new_n348_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(KEYINPUT94), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n346_), .ZN(new_n359_));
  AND4_X1   g158(.A1(KEYINPUT94), .A2(new_n343_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n354_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n302_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n354_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n341_), .B1(KEYINPUT94), .B2(new_n355_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n365_), .B2(new_n360_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n299_), .A2(new_n301_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n356_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n270_), .B1(new_n363_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n325_), .A2(new_n328_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n313_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT4), .B1(new_n371_), .B2(new_n297_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n297_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n329_), .A2(new_n296_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n372_), .B1(new_n375_), .B2(KEYINPUT4), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT99), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n375_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n377_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT99), .ZN(new_n381_));
  INV_X1    g180(.A(new_n377_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n381_), .B(new_n382_), .C1(new_n384_), .C2(new_n372_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n378_), .A2(new_n380_), .A3(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT0), .B(G57gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G85gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(G1gat), .B(G29gat), .Z(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(new_n389_), .Z(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n390_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n378_), .A2(new_n392_), .A3(new_n380_), .A4(new_n385_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n379_), .A2(new_n382_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n396_), .B(new_n390_), .C1(new_n376_), .C2(new_n382_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n261_), .B1(new_n398_), .B2(KEYINPUT33), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n393_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT32), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n260_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n266_), .A2(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n405_), .B(KEYINPUT100), .Z(new_n406_));
  OAI211_X1 g205(.A(new_n394_), .B(new_n406_), .C1(new_n256_), .C2(new_n404_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n367_), .B1(new_n402_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n357_), .A2(new_n362_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n369_), .A2(new_n395_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G229gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G29gat), .B(G36gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(new_n276_), .ZN(new_n413_));
  INV_X1    g212(.A(G50gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G15gat), .B(G22gat), .ZN(new_n416_));
  INV_X1    g215(.A(G1gat), .ZN(new_n417_));
  INV_X1    g216(.A(G8gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT14), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G1gat), .B(G8gat), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(new_n421_), .Z(new_n422_));
  NAND2_X1  g221(.A1(new_n415_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n415_), .A2(KEYINPUT15), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n413_), .B(G50gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT15), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n411_), .B(new_n423_), .C1(new_n428_), .C2(new_n422_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n422_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n423_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n411_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G113gat), .B(G141gat), .ZN(new_n436_));
  INV_X1    g235(.A(G169gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G197gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT81), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT82), .Z(new_n442_));
  XNOR2_X1  g241(.A(new_n435_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n410_), .A2(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n445_), .A2(KEYINPUT102), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(KEYINPUT102), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G99gat), .A2(G106gat), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT64), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n452_), .B1(new_n456_), .B2(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G85gat), .B(G92gat), .Z(new_n463_));
  INV_X1    g262(.A(KEYINPUT8), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT65), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT7), .ZN(new_n468_));
  INV_X1    g267(.A(G99gat), .ZN(new_n469_));
  INV_X1    g268(.A(G106gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n449_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n455_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n459_), .A2(KEYINPUT64), .A3(new_n460_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT65), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n465_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n467_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT66), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n459_), .A2(KEYINPUT66), .A3(new_n460_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n452_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n463_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT8), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT67), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n483_), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n478_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT11), .ZN(new_n489_));
  OR2_X1    g288(.A1(G57gat), .A2(G64gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G57gat), .A2(G64gat), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n493_), .A2(new_n494_), .A3(G78gat), .ZN(new_n495_));
  INV_X1    g294(.A(G78gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT68), .ZN(new_n497_));
  INV_X1    g296(.A(G71gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n496_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n492_), .B1(new_n495_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n491_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(G57gat), .A2(G64gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT11), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n490_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n506_));
  OAI21_X1  g305(.A(G78gat), .B1(new_n493_), .B2(new_n494_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n499_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n502_), .A2(new_n509_), .A3(KEYINPUT69), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT69), .B1(new_n502_), .B2(new_n509_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n463_), .A2(KEYINPUT9), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT10), .B(G99gat), .ZN(new_n516_));
  OAI221_X1 g315(.A(new_n514_), .B1(KEYINPUT9), .B2(new_n515_), .C1(G106gat), .C2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n456_), .A2(new_n461_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n488_), .A2(new_n513_), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT67), .B1(new_n483_), .B2(KEYINPUT8), .ZN(new_n524_));
  AOI211_X1 g323(.A(new_n485_), .B(new_n464_), .C1(new_n482_), .C2(new_n463_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n519_), .B1(new_n526_), .B2(new_n478_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT71), .B1(new_n527_), .B2(new_n513_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n488_), .A2(new_n520_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n512_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(KEYINPUT70), .A3(new_n513_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n523_), .A2(new_n528_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G230gat), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(new_n334_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT72), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT74), .B(KEYINPUT12), .Z(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n527_), .B2(new_n513_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n502_), .A2(new_n509_), .A3(KEYINPUT12), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT73), .B1(new_n527_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT73), .ZN(new_n542_));
  INV_X1    g341(.A(new_n540_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n529_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  AND4_X1   g343(.A1(new_n521_), .A2(new_n539_), .A3(new_n541_), .A4(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n535_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n533_), .A2(new_n548_), .A3(new_n535_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n537_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G120gat), .B(G148gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(new_n232_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT5), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n223_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n537_), .A2(new_n547_), .A3(new_n549_), .A4(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT13), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(KEYINPUT75), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n559_), .A2(KEYINPUT75), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n558_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT76), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n424_), .A2(new_n427_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n529_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT78), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT34), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(KEYINPUT35), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n527_), .B2(new_n415_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT79), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(KEYINPUT35), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT77), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(G134gat), .ZN(new_n581_));
  INV_X1    g380(.A(G162gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT36), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n574_), .A2(new_n578_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n579_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n579_), .B2(new_n586_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT37), .B1(new_n587_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n579_), .A2(new_n586_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n589_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n579_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n592_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n422_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT80), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n513_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT16), .B(G183gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(G211gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT17), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n502_), .A2(new_n509_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n600_), .B(new_n609_), .Z(new_n610_));
  INV_X1    g409(.A(KEYINPUT17), .ZN(new_n611_));
  OR3_X1    g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n606_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n598_), .A2(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n448_), .A2(new_n565_), .A3(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n417_), .A3(new_n394_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT38), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n587_), .A2(new_n591_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT103), .ZN(new_n619_));
  INV_X1    g418(.A(new_n613_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n445_), .A2(new_n564_), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n395_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n617_), .A2(new_n623_), .ZN(G1324gat));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n625_));
  INV_X1    g424(.A(new_n270_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(G8gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n628_), .B1(new_n627_), .B2(G8gat), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n625_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(G8gat), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT104), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(KEYINPUT39), .A3(new_n629_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n615_), .A2(new_n418_), .A3(new_n270_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n632_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n632_), .A2(new_n635_), .A3(KEYINPUT40), .A4(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1325gat));
  OAI21_X1  g440(.A(G15gat), .B1(new_n622_), .B2(new_n302_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT41), .Z(new_n643_));
  INV_X1    g442(.A(G15gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n615_), .A2(new_n644_), .A3(new_n367_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT105), .ZN(G1326gat));
  INV_X1    g446(.A(G22gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n409_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n615_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G22gat), .B1(new_n622_), .B2(new_n409_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(G1327gat));
  AND3_X1   g454(.A1(new_n366_), .A2(new_n367_), .A3(new_n356_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n367_), .B1(new_n366_), .B2(new_n356_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n395_), .B(new_n626_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n402_), .A2(new_n407_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n302_), .A3(new_n409_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n598_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n592_), .A2(new_n597_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT43), .B1(new_n667_), .B2(KEYINPUT107), .ZN(new_n668_));
  INV_X1    g467(.A(new_n564_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n444_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n665_), .A2(new_n668_), .A3(new_n613_), .A4(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n672_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n394_), .A3(new_n674_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(KEYINPUT108), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(KEYINPUT108), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(G29gat), .A3(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n619_), .A2(new_n620_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n448_), .A2(new_n564_), .A3(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n395_), .A2(G29gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT109), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n680_), .B2(new_n682_), .ZN(G1328gat));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n626_), .A2(G36gat), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n680_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n679_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n689_), .A2(KEYINPUT45), .A3(new_n564_), .A4(new_n685_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n673_), .A2(new_n270_), .A3(new_n674_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n691_), .B(KEYINPUT46), .C1(new_n692_), .C2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n693_), .A2(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n687_), .A2(new_n690_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n695_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n698_), .ZN(G1329gat));
  NAND4_X1  g498(.A1(new_n689_), .A2(new_n276_), .A3(new_n564_), .A4(new_n367_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n673_), .A2(new_n367_), .A3(new_n674_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n276_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n700_), .B(KEYINPUT47), .C1(new_n701_), .C2(new_n276_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1330gat));
  OAI21_X1  g505(.A(new_n414_), .B1(new_n680_), .B2(new_n409_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n673_), .A2(G50gat), .A3(new_n649_), .A4(new_n674_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT110), .ZN(G1331gat));
  NAND3_X1  g509(.A1(new_n666_), .A2(new_n620_), .A3(new_n444_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n410_), .A2(new_n711_), .A3(new_n564_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G57gat), .B1(new_n712_), .B2(new_n394_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n565_), .A2(new_n443_), .A3(new_n410_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(new_n621_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(new_n394_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n713_), .B1(new_n716_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g516(.A(G64gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n715_), .B2(new_n270_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT48), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n712_), .A2(new_n718_), .A3(new_n270_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1333gat));
  AOI21_X1  g521(.A(new_n498_), .B1(new_n715_), .B2(new_n367_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT49), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n712_), .A2(new_n498_), .A3(new_n367_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1334gat));
  AOI21_X1  g525(.A(new_n496_), .B1(new_n715_), .B2(new_n649_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT50), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n712_), .A2(new_n496_), .A3(new_n649_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1335gat));
  AND2_X1   g529(.A1(new_n714_), .A2(new_n679_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n394_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n664_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n667_), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT111), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n665_), .A2(new_n736_), .A3(new_n668_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n669_), .A2(new_n613_), .A3(new_n444_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT112), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n394_), .A2(G85gat), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT113), .Z(new_n744_));
  AOI21_X1  g543(.A(new_n732_), .B1(new_n742_), .B2(new_n744_), .ZN(G1336gat));
  AOI21_X1  g544(.A(G92gat), .B1(new_n731_), .B2(new_n270_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n741_), .A2(new_n626_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(G92gat), .ZN(G1337gat));
  NAND4_X1  g547(.A1(new_n735_), .A2(new_n367_), .A3(new_n740_), .A4(new_n737_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G99gat), .ZN(new_n750_));
  INV_X1    g549(.A(new_n516_), .ZN(new_n751_));
  AND4_X1   g550(.A1(new_n751_), .A2(new_n714_), .A3(new_n367_), .A4(new_n679_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n750_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT114), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n750_), .A2(new_n756_), .A3(new_n753_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT51), .B1(new_n755_), .B2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT114), .B(new_n752_), .C1(new_n749_), .C2(G99gat), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n758_), .A2(new_n762_), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n731_), .A2(new_n470_), .A3(new_n649_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n740_), .A2(new_n649_), .A3(new_n668_), .A4(new_n665_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G106gat), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g569(.A1(new_n711_), .A2(KEYINPUT54), .A3(new_n669_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n598_), .A2(new_n613_), .A3(new_n443_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(new_n564_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n771_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n542_), .B1(new_n529_), .B2(new_n543_), .ZN(new_n776_));
  AOI211_X1 g575(.A(KEYINPUT73), .B(new_n540_), .C1(new_n488_), .C2(new_n520_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n519_), .B(new_n512_), .C1(new_n526_), .C2(new_n478_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n529_), .A2(new_n512_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(new_n538_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n778_), .A2(KEYINPUT55), .A3(new_n781_), .A4(new_n546_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n545_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n546_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n539_), .A2(new_n541_), .A3(new_n544_), .A4(new_n521_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n535_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n535_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n555_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n784_), .B(new_n785_), .C1(new_n790_), .C2(new_n789_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n555_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n557_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n555_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(KEYINPUT116), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n801_), .A3(new_n443_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n422_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n423_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n803_), .A2(new_n411_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n432_), .A2(new_n411_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n440_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n440_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n803_), .A2(new_n433_), .A3(new_n804_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n434_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n809_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n808_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n808_), .B2(new_n812_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT118), .B1(new_n558_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n819_), .B(new_n816_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n802_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n619_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n822_), .B(new_n619_), .C1(new_n824_), .C2(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n794_), .A2(new_n797_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n817_), .B2(new_n557_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n799_), .A2(KEYINPUT120), .A3(new_n816_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n828_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(KEYINPUT121), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(KEYINPUT121), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n828_), .B(new_n835_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n836_), .A3(new_n598_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n826_), .A2(new_n827_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n775_), .B1(new_n838_), .B2(new_n613_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n270_), .A2(new_n395_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n839_), .A2(new_n368_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n443_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT122), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n838_), .A2(new_n613_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n775_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n841_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n847_), .B1(new_n850_), .B2(new_n656_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NOR4_X1   g652(.A1(new_n839_), .A2(new_n368_), .A3(new_n841_), .A4(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n845_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n848_), .A2(new_n849_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n856_), .A2(new_n656_), .A3(new_n840_), .A4(new_n852_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(KEYINPUT123), .C1(new_n842_), .C2(new_n847_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n444_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n844_), .B1(new_n859_), .B2(new_n843_), .ZN(G1340gat));
  NOR2_X1   g659(.A1(new_n851_), .A2(new_n854_), .ZN(new_n861_));
  OAI21_X1  g660(.A(G120gat), .B1(new_n861_), .B2(new_n565_), .ZN(new_n862_));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n564_), .B2(KEYINPUT60), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n842_), .B(new_n864_), .C1(KEYINPUT60), .C2(new_n863_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1341gat));
  INV_X1    g665(.A(G127gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n842_), .A2(new_n867_), .A3(new_n620_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n613_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1342gat));
  NOR2_X1   g669(.A1(new_n619_), .A2(G134gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n842_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n666_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n873_));
  INV_X1    g672(.A(G134gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(G1343gat));
  NAND2_X1  g674(.A1(new_n850_), .A2(new_n657_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n444_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n309_), .ZN(G1344gat));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n565_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n310_), .ZN(G1345gat));
  NOR2_X1   g679(.A1(new_n876_), .A2(new_n613_), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT61), .B(G155gat), .Z(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  NOR3_X1   g682(.A1(new_n876_), .A2(new_n582_), .A3(new_n666_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n876_), .A2(new_n619_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n582_), .B2(new_n885_), .ZN(G1347gat));
  NOR3_X1   g685(.A1(new_n839_), .A2(new_n394_), .A3(new_n626_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n656_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G169gat), .B1(new_n888_), .B2(new_n444_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n888_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n443_), .A3(new_n222_), .ZN(new_n893_));
  OAI211_X1 g692(.A(KEYINPUT62), .B(G169gat), .C1(new_n888_), .C2(new_n444_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n891_), .A2(new_n893_), .A3(new_n894_), .ZN(G1348gat));
  AOI21_X1  g694(.A(G176gat), .B1(new_n892_), .B2(new_n669_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n887_), .A2(G176gat), .A3(new_n656_), .ZN(new_n897_));
  OR3_X1    g696(.A1(new_n897_), .A2(KEYINPUT124), .A3(new_n565_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT124), .B1(new_n897_), .B2(new_n565_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n896_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  NOR2_X1   g699(.A1(new_n888_), .A2(new_n613_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n202_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n211_), .B2(new_n901_), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n888_), .B2(new_n666_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n203_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n619_), .A2(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT125), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n904_), .B1(new_n888_), .B2(new_n907_), .ZN(G1351gat));
  NAND2_X1  g707(.A1(new_n887_), .A2(new_n657_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n444_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n439_), .ZN(G1352gat));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n565_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n232_), .ZN(G1353gat));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914_));
  NAND2_X1  g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n620_), .A2(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n887_), .B(new_n657_), .C1(new_n914_), .C2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n914_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921_));
  NOR2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n921_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n924_), .B(new_n925_), .C1(new_n917_), .C2(new_n919_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n923_), .A2(new_n926_), .ZN(G1354gat));
  NOR2_X1   g726(.A1(new_n909_), .A2(new_n619_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(G218gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n909_), .A2(new_n666_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(G218gat), .B2(new_n930_), .ZN(G1355gat));
endmodule


