//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n963_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G85gat), .B(G92gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n207_), .B(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT64), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n208_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT7), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n213_), .B1(new_n221_), .B2(new_n205_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n205_), .A2(new_n213_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n208_), .B2(new_n220_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n212_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G29gat), .B(G36gat), .Z(new_n226_));
  XOR2_X1   g025(.A(G43gat), .B(G50gat), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G29gat), .B(G36gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT15), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n225_), .A2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n232_), .B(new_n212_), .C1(new_n222_), .C2(new_n224_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G232gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT34), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT35), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n238_), .A2(new_n239_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT69), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n234_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n241_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n234_), .B1(new_n245_), .B2(KEYINPUT67), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(KEYINPUT67), .B2(new_n245_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n244_), .B1(new_n247_), .B2(new_n242_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G190gat), .B(G218gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT68), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G134gat), .B(G162gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(KEYINPUT36), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n252_), .B(KEYINPUT36), .Z(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT70), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n248_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT37), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n257_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n247_), .A2(new_n242_), .ZN(new_n262_));
  OAI211_X1 g061(.A(KEYINPUT71), .B(new_n261_), .C1(new_n262_), .C2(new_n244_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n263_), .A2(new_n254_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT37), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(new_n248_), .B2(new_n257_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n264_), .A2(KEYINPUT72), .A3(new_n265_), .A4(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n263_), .A2(new_n267_), .A3(new_n254_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(KEYINPUT37), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n260_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT75), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G1gat), .B(G8gat), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT73), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT73), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G15gat), .B(G22gat), .ZN(new_n278_));
  INV_X1    g077(.A(G1gat), .ZN(new_n279_));
  INV_X1    g078(.A(G8gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT14), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n275_), .A2(new_n281_), .A3(new_n278_), .A4(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G57gat), .B(G64gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT11), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT65), .B(G71gat), .ZN(new_n290_));
  INV_X1    g089(.A(G78gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n293_), .B1(new_n294_), .B2(new_n292_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n287_), .B(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G127gat), .B(G155gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(G183gat), .B(G211gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT17), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n296_), .A2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n301_), .A2(KEYINPUT17), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n273_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n305_), .A2(new_n273_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n272_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G230gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n225_), .A2(new_n295_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n313_), .A2(KEYINPUT12), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n292_), .A2(new_n294_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n315_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n316_), .B(new_n212_), .C1(new_n222_), .C2(new_n224_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n317_), .A3(KEYINPUT12), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n312_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n311_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G120gat), .B(G148gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G176gat), .B(G204gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n321_), .A2(new_n326_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT13), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(KEYINPUT13), .A3(new_n328_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n310_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT76), .ZN(new_n335_));
  OR3_X1    g134(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n336_));
  INV_X1    g135(.A(G169gat), .ZN(new_n337_));
  INV_X1    g136(.A(G176gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n336_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(G183gat), .A3(G190gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT85), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n342_), .A2(KEYINPUT85), .A3(G183gat), .A4(G190gat), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT84), .B1(new_n348_), .B2(KEYINPUT23), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n341_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n354_));
  INV_X1    g153(.A(G183gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(KEYINPUT25), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT81), .B1(new_n357_), .B2(G183gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(G183gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G190gat), .ZN(new_n361_));
  AND4_X1   g160(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .A4(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT82), .B(G190gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(KEYINPUT26), .ZN(new_n365_));
  INV_X1    g164(.A(G190gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT82), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G190gat), .ZN(new_n369_));
  AND4_X1   g168(.A1(new_n363_), .A2(new_n367_), .A3(new_n369_), .A4(KEYINPUT26), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n362_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n337_), .A2(KEYINPUT22), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT22), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G169gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n374_), .A3(new_n338_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n339_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n348_), .A2(KEYINPUT23), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n343_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n367_), .A2(new_n369_), .A3(new_n355_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n377_), .A2(KEYINPUT86), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n375_), .A2(new_n382_), .A3(new_n376_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n353_), .A2(new_n371_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G71gat), .B(G99gat), .ZN(new_n385_));
  INV_X1    g184(.A(G43gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n384_), .B(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G127gat), .B(G134gat), .Z(new_n389_));
  XOR2_X1   g188(.A(G113gat), .B(G120gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n388_), .B(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(G15gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT30), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT31), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n392_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n392_), .A2(new_n398_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT27), .ZN(new_n403_));
  XOR2_X1   g202(.A(G8gat), .B(G36gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G197gat), .A2(G204gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT89), .B(G197gat), .ZN(new_n411_));
  INV_X1    g210(.A(G204gat), .ZN(new_n412_));
  OAI211_X1 g211(.A(KEYINPUT91), .B(new_n410_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G211gat), .B(G218gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT21), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G197gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT89), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT89), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G197gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G204gat), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT91), .B1(new_n423_), .B2(new_n410_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT92), .B1(new_n417_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT91), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n412_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n409_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT92), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n413_), .A4(new_n416_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT21), .B1(new_n423_), .B2(new_n410_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n419_), .A2(new_n421_), .A3(new_n412_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n415_), .B1(G197gat), .B2(G204gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n414_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT90), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n415_), .B1(new_n427_), .B2(new_n409_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n414_), .A4(new_n435_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n384_), .B1(new_n431_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT19), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n442_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n425_), .A2(new_n430_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n339_), .A2(new_n340_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT25), .B(G183gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT26), .B(G190gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n448_), .A2(new_n451_), .A3(new_n379_), .A4(new_n336_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT93), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n348_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n345_), .B(new_n346_), .C1(new_n455_), .C2(new_n349_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n355_), .A2(new_n366_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT95), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n456_), .A2(KEYINPUT95), .A3(new_n457_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n339_), .A2(KEYINPUT94), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n339_), .A2(KEYINPUT94), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n372_), .A2(new_n374_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n463_), .A2(new_n464_), .B1(new_n465_), .B2(new_n338_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT96), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n456_), .A2(KEYINPUT95), .A3(new_n457_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT95), .B1(new_n456_), .B2(new_n457_), .ZN(new_n469_));
  OAI211_X1 g268(.A(KEYINPUT96), .B(new_n466_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n447_), .B(new_n454_), .C1(new_n467_), .C2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n443_), .B1(new_n447_), .B2(new_n384_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n466_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n453_), .B1(new_n476_), .B2(new_n470_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n473_), .B1(new_n477_), .B2(new_n447_), .ZN(new_n478_));
  AOI221_X4 g277(.A(new_n408_), .B1(new_n446_), .B2(new_n472_), .C1(new_n478_), .C2(new_n445_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n408_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n445_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n446_), .A2(new_n472_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n403_), .B1(new_n479_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G1gat), .B(G29gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G85gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT0), .B(G57gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G225gat), .A2(G233gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT98), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G155gat), .A2(G162gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G155gat), .A2(G162gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT87), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(G155gat), .A3(G162gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n493_), .B1(new_n498_), .B2(KEYINPUT1), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT1), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G141gat), .A2(G148gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G141gat), .A2(G148gat), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT2), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n503_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n509_), .A2(new_n511_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n493_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT88), .B1(new_n498_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n517_));
  AOI211_X1 g316(.A(new_n517_), .B(new_n493_), .C1(new_n495_), .C2(new_n497_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n514_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n391_), .B1(new_n507_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT4), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n492_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n391_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n514_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n498_), .A2(new_n515_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n517_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n498_), .A2(KEYINPUT88), .A3(new_n515_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n524_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n506_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n523_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n507_), .A2(new_n519_), .A3(new_n391_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT4), .A3(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n522_), .A2(new_n533_), .A3(KEYINPUT99), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n531_), .A2(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n490_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT99), .B1(new_n522_), .B2(new_n533_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n489_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n522_), .A2(new_n533_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT99), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n542_), .A2(new_n488_), .A3(new_n536_), .A4(new_n534_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n539_), .A2(KEYINPUT103), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT103), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n545_), .B(new_n489_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n481_), .A2(new_n480_), .A3(new_n482_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n445_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n431_), .A2(new_n441_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n384_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n443_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n447_), .A2(new_n452_), .A3(new_n474_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n549_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT20), .B1(new_n550_), .B2(new_n551_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n454_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n556_), .B2(new_n550_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n554_), .B1(new_n557_), .B2(new_n549_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n548_), .B(KEYINPUT27), .C1(new_n558_), .C2(new_n480_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n484_), .A2(new_n547_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n507_), .A2(new_n519_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n561_), .A2(KEYINPUT29), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT28), .Z(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(KEYINPUT29), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n550_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n562_), .B(KEYINPUT28), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(new_n550_), .A3(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G228gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(new_n291_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n203_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G22gat), .B(G50gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n566_), .A2(new_n568_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n402_), .B1(new_n560_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT100), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(KEYINPUT33), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n543_), .A2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n534_), .A2(new_n536_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n582_), .A2(new_n488_), .A3(new_n542_), .A4(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n481_), .A2(new_n482_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n408_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n535_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n492_), .B1(new_n587_), .B2(KEYINPUT101), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(KEYINPUT101), .B2(new_n587_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n533_), .B(new_n490_), .C1(KEYINPUT4), .C2(new_n531_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n489_), .A3(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n584_), .A2(new_n586_), .A3(new_n548_), .A4(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n574_), .A2(new_n575_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT102), .B1(new_n558_), .B2(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n447_), .A2(new_n452_), .A3(new_n474_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT20), .B1(new_n447_), .B2(new_n384_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n445_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n478_), .B2(new_n445_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT102), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(KEYINPUT32), .A4(new_n480_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n481_), .A2(new_n594_), .A3(new_n482_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n595_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n592_), .B(new_n593_), .C1(new_n603_), .C2(new_n547_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n577_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT104), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT104), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n577_), .A2(new_n607_), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n484_), .A2(new_n559_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n576_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n547_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n401_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n606_), .A2(new_n608_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n283_), .A2(new_n284_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n232_), .B(KEYINPUT77), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT77), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n232_), .B(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n285_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G229gat), .A2(G233gat), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT78), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n614_), .A2(new_n233_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT79), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G113gat), .B(G141gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G169gat), .B(G197gat), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n628_), .B(new_n629_), .Z(new_n630_));
  NOR2_X1   g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n624_), .A2(new_n626_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT79), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n634_), .A3(new_n630_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(KEYINPUT80), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT80), .ZN(new_n637_));
  INV_X1    g436(.A(new_n635_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(new_n631_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n613_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT76), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n310_), .A2(new_n643_), .A3(new_n333_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n335_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n645_), .A2(G1gat), .A3(new_n547_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(KEYINPUT38), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT107), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n638_), .A2(new_n631_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n333_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(new_n309_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n270_), .A2(KEYINPUT105), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n263_), .A2(new_n267_), .A3(new_n654_), .A4(new_n254_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT106), .B1(new_n613_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n610_), .A2(new_n612_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n560_), .A2(new_n576_), .ZN(new_n660_));
  AND4_X1   g459(.A1(new_n607_), .A2(new_n660_), .A3(new_n604_), .A4(new_n401_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n607_), .B1(new_n577_), .B2(new_n604_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n664_), .A3(new_n656_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n652_), .B1(new_n658_), .B2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n279_), .B1(new_n666_), .B2(new_n611_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n646_), .B2(KEYINPUT38), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n648_), .A2(new_n668_), .ZN(G1324gat));
  INV_X1    g468(.A(KEYINPUT109), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n280_), .B1(new_n666_), .B2(new_n609_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT39), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT110), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n674_), .A3(new_n672_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n665_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n664_), .B1(new_n663_), .B2(new_n656_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n609_), .B(new_n651_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G8gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(KEYINPUT109), .A3(KEYINPUT39), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n672_), .A3(G8gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT110), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n673_), .A2(new_n675_), .A3(new_n680_), .A4(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n609_), .A2(new_n280_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n645_), .A2(KEYINPUT108), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT108), .B1(new_n645_), .B2(new_n684_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n683_), .A2(KEYINPUT40), .A3(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1325gat));
  AOI21_X1  g491(.A(new_n394_), .B1(new_n666_), .B2(new_n402_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(KEYINPUT41), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(KEYINPUT41), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n402_), .A2(new_n394_), .ZN(new_n696_));
  OAI22_X1  g495(.A1(new_n694_), .A2(new_n695_), .B1(new_n645_), .B2(new_n696_), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n666_), .A2(new_n576_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G22gat), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT42), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(KEYINPUT42), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n593_), .A2(G22gat), .ZN(new_n702_));
  OAI22_X1  g501(.A1(new_n700_), .A2(new_n701_), .B1(new_n645_), .B2(new_n702_), .ZN(G1327gat));
  NOR2_X1   g502(.A1(new_n656_), .A2(new_n308_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n642_), .A2(new_n333_), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n611_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n663_), .A2(new_n707_), .A3(new_n272_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n663_), .A2(KEYINPUT111), .A3(new_n707_), .A4(new_n272_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n268_), .A2(new_n271_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n259_), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT43), .B1(new_n613_), .B2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n710_), .A2(new_n711_), .A3(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n650_), .A2(new_n308_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n715_), .A2(KEYINPUT44), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT44), .B1(new_n715_), .B2(new_n716_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n611_), .A2(G29gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n706_), .B1(new_n719_), .B2(new_n720_), .ZN(G1328gat));
  INV_X1    g520(.A(new_n609_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(G36gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n705_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n705_), .A2(KEYINPUT45), .A3(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n717_), .A2(new_n718_), .A3(new_n722_), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(KEYINPUT112), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n733_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n715_), .A2(new_n716_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n715_), .A2(KEYINPUT44), .A3(new_n716_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n609_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n728_), .B1(new_n740_), .B2(G36gat), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n735_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n734_), .A2(new_n743_), .ZN(G1329gat));
  AOI21_X1  g543(.A(G43gat), .B1(new_n705_), .B2(new_n402_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n401_), .A2(new_n386_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n719_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(G1330gat));
  NOR2_X1   g548(.A1(new_n593_), .A2(G50gat), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n705_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n738_), .A2(new_n576_), .A3(new_n739_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(G50gat), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT114), .ZN(G1331gat));
  NAND3_X1  g553(.A1(new_n636_), .A2(new_n308_), .A3(new_n639_), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n333_), .B(new_n755_), .C1(new_n658_), .C2(new_n665_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G57gat), .B1(new_n757_), .B2(new_n547_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n613_), .A2(new_n333_), .A3(new_n649_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(new_n310_), .ZN(new_n760_));
  INV_X1    g559(.A(G57gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n611_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(new_n762_), .ZN(G1332gat));
  INV_X1    g562(.A(G64gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n764_), .A3(new_n609_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G64gat), .B1(new_n757_), .B2(new_n722_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT48), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT48), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n765_), .B1(new_n767_), .B2(new_n768_), .ZN(G1333gat));
  INV_X1    g568(.A(G71gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n760_), .A2(new_n770_), .A3(new_n402_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n756_), .A2(new_n402_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(G71gat), .ZN(new_n774_));
  AOI211_X1 g573(.A(KEYINPUT49), .B(new_n770_), .C1(new_n756_), .C2(new_n402_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT115), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n771_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1334gat));
  NAND3_X1  g579(.A1(new_n760_), .A2(new_n291_), .A3(new_n576_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G78gat), .B1(new_n757_), .B2(new_n593_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(KEYINPUT50), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(KEYINPUT50), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n783_), .B2(new_n784_), .ZN(G1335gat));
  AND2_X1   g584(.A1(new_n759_), .A2(new_n704_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n209_), .A3(new_n611_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n333_), .A2(new_n308_), .A3(new_n649_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n715_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n715_), .A2(KEYINPUT116), .A3(new_n788_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n547_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n787_), .B1(new_n793_), .B2(new_n209_), .ZN(G1336gat));
  NAND3_X1  g593(.A1(new_n786_), .A2(new_n210_), .A3(new_n609_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n722_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n210_), .ZN(G1337gat));
  NAND3_X1  g596(.A1(new_n786_), .A2(new_n202_), .A3(new_n402_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n401_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n799_));
  INV_X1    g598(.A(G99gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT51), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n798_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1338gat));
  NAND3_X1  g604(.A1(new_n786_), .A2(new_n203_), .A3(new_n576_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n715_), .A2(new_n576_), .A3(new_n788_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n807_), .A2(G106gat), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n807_), .B2(G106gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g611(.A1(new_n609_), .A2(new_n576_), .A3(new_n401_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n620_), .A2(new_n621_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n625_), .A2(new_n619_), .A3(new_n622_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  MUX2_X1   g615(.A(new_n816_), .B(new_n633_), .S(new_n630_), .Z(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n327_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n314_), .A2(new_n312_), .A3(new_n318_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT55), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(new_n319_), .ZN(new_n821_));
  AOI211_X1 g620(.A(KEYINPUT55), .B(new_n312_), .C1(new_n314_), .C2(new_n318_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT119), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n314_), .A2(new_n318_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n311_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT55), .A3(new_n819_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n822_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n823_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT56), .B1(new_n830_), .B2(new_n326_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n818_), .B1(new_n831_), .B2(KEYINPUT120), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n821_), .A2(KEYINPUT119), .A3(new_n822_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n828_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n326_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n326_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n832_), .A2(new_n840_), .A3(KEYINPUT58), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n832_), .A2(new_n840_), .A3(KEYINPUT121), .A4(KEYINPUT58), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT58), .B1(new_n832_), .B2(new_n840_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n713_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n649_), .A2(new_n327_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n329_), .A2(new_n817_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n656_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n656_), .B(KEYINPUT57), .C1(new_n850_), .C2(new_n852_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n308_), .B1(new_n848_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n755_), .A2(KEYINPUT118), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n636_), .A2(new_n639_), .A3(new_n861_), .A4(new_n308_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n333_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n859_), .B1(new_n864_), .B2(new_n713_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n863_), .A2(new_n272_), .A3(KEYINPUT54), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n611_), .B(new_n813_), .C1(new_n858_), .C2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(G113gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n649_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n868_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n855_), .A2(new_n856_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n875_));
  OAI22_X1  g674(.A1(new_n875_), .A2(new_n308_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n876_), .A2(KEYINPUT59), .A3(new_n611_), .A4(new_n813_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n641_), .B1(new_n873_), .B2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n871_), .B1(new_n878_), .B2(new_n870_), .ZN(G1340gat));
  AOI21_X1  g678(.A(new_n333_), .B1(new_n873_), .B2(new_n877_), .ZN(new_n880_));
  INV_X1    g679(.A(G120gat), .ZN(new_n881_));
  INV_X1    g680(.A(new_n333_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n883_));
  AOI21_X1  g682(.A(G120gat), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n883_), .B2(G120gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT122), .B1(new_n869_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887_));
  INV_X1    g686(.A(new_n885_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n868_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  OAI22_X1  g688(.A1(new_n880_), .A2(new_n881_), .B1(new_n886_), .B2(new_n889_), .ZN(G1341gat));
  INV_X1    g689(.A(G127gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n869_), .A2(new_n891_), .A3(new_n308_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n309_), .B1(new_n873_), .B2(new_n877_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1342gat));
  AOI21_X1  g693(.A(G134gat), .B1(new_n869_), .B2(new_n657_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n873_), .A2(new_n877_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n272_), .A2(G134gat), .ZN(new_n897_));
  XOR2_X1   g696(.A(new_n897_), .B(KEYINPUT123), .Z(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n896_), .B2(new_n898_), .ZN(G1343gat));
  NOR2_X1   g698(.A1(new_n593_), .A2(new_n402_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n609_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n876_), .A2(new_n611_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n649_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT124), .B(G141gat), .Z(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1344gat));
  NOR2_X1   g706(.A1(new_n903_), .A2(new_n333_), .ZN(new_n908_));
  INV_X1    g707(.A(G148gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1345gat));
  NOR2_X1   g709(.A1(new_n903_), .A2(new_n309_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT61), .B(G155gat), .Z(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n903_), .B2(new_n713_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n656_), .A2(G162gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n903_), .B2(new_n915_), .ZN(G1347gat));
  NAND3_X1  g715(.A1(new_n612_), .A2(new_n593_), .A3(new_n609_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n876_), .A2(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919_), .B2(new_n904_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n921_), .ZN(new_n923_));
  OAI211_X1 g722(.A(G169gat), .B(new_n923_), .C1(new_n919_), .C2(new_n904_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n876_), .A2(new_n465_), .A3(new_n649_), .A4(new_n918_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n922_), .A2(new_n924_), .A3(new_n925_), .ZN(G1348gat));
  NAND3_X1  g725(.A1(new_n876_), .A2(new_n882_), .A3(new_n918_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g727(.A1(new_n876_), .A2(new_n308_), .A3(new_n918_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(new_n449_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n355_), .B2(new_n929_), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n919_), .B2(new_n713_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n657_), .A2(new_n450_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n919_), .B2(new_n933_), .ZN(G1351gat));
  NAND2_X1  g733(.A1(new_n848_), .A2(new_n857_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n867_), .B1(new_n935_), .B2(new_n309_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n901_), .A2(new_n611_), .A3(new_n722_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(KEYINPUT126), .B1(new_n936_), .B2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n940_), .B(new_n937_), .C1(new_n858_), .C2(new_n867_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942_), .B2(new_n649_), .ZN(new_n943_));
  AOI211_X1 g742(.A(new_n418_), .B(new_n904_), .C1(new_n939_), .C2(new_n941_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1352gat));
  AOI21_X1  g744(.A(new_n940_), .B1(new_n876_), .B2(new_n937_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n941_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n882_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(G204gat), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n942_), .A2(new_n412_), .A3(new_n882_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1353gat));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  AND2_X1   g753(.A1(new_n308_), .A2(new_n954_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n953_), .B1(new_n942_), .B2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n955_), .ZN(new_n957_));
  AOI211_X1 g756(.A(new_n952_), .B(new_n957_), .C1(new_n939_), .C2(new_n941_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n956_), .A2(new_n958_), .ZN(G1354gat));
  NAND2_X1  g758(.A1(new_n942_), .A2(new_n657_), .ZN(new_n960_));
  INV_X1    g759(.A(G218gat), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n272_), .A2(G218gat), .ZN(new_n962_));
  XOR2_X1   g761(.A(new_n962_), .B(KEYINPUT127), .Z(new_n963_));
  AOI22_X1  g762(.A1(new_n960_), .A2(new_n961_), .B1(new_n942_), .B2(new_n963_), .ZN(G1355gat));
endmodule


