//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G78gat), .Z(new_n204_));
  OR2_X1    g003(.A1(G57gat), .A2(G64gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G57gat), .A2(G64gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n203_), .B1(new_n204_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n206_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n204_), .A2(new_n208_), .A3(new_n203_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n211_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n212_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(new_n209_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n221_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT8), .B1(new_n227_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT10), .B(G99gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT64), .B1(new_n232_), .B2(G106gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n224_), .A2(KEYINPUT10), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT10), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G99gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n225_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n233_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n228_), .A2(KEYINPUT9), .A3(new_n229_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n229_), .A2(KEYINPUT9), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n221_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT65), .B1(new_n240_), .B2(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n221_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n233_), .A4(new_n239_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n231_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n226_), .A2(new_n222_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT66), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n226_), .A2(new_n251_), .A3(new_n222_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n221_), .A3(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(KEYINPUT8), .A3(new_n230_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n248_), .A2(KEYINPUT68), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT68), .B1(new_n248_), .B2(new_n254_), .ZN(new_n256_));
  OAI211_X1 g055(.A(KEYINPUT12), .B(new_n218_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n231_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n238_), .B1(new_n237_), .B2(new_n225_), .ZN(new_n259_));
  AOI211_X1 g058(.A(KEYINPUT64), .B(G106gat), .C1(new_n234_), .C2(new_n236_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n246_), .B1(new_n261_), .B2(new_n245_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n240_), .A2(KEYINPUT65), .A3(new_n243_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n258_), .B(new_n254_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT12), .B1(new_n264_), .B2(new_n218_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n218_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n257_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n268_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n217_), .B1(new_n248_), .B2(new_n254_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n270_), .B1(new_n266_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT5), .B(G176gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G204gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G120gat), .B(G148gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  OAI21_X1  g076(.A(new_n202_), .B1(new_n273_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n269_), .A2(KEYINPUT69), .A3(new_n272_), .A4(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n273_), .A2(new_n277_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT13), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n286_));
  INV_X1    g085(.A(G29gat), .ZN(new_n287_));
  INV_X1    g086(.A(G36gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G29gat), .A2(G36gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G50gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G43gat), .ZN(new_n293_));
  INV_X1    g092(.A(G43gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(G50gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n293_), .A2(new_n295_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n299_), .A3(KEYINPUT15), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT15), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n296_), .A2(new_n291_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(new_n298_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT14), .ZN(new_n305_));
  INV_X1    g104(.A(G8gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT73), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G8gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n305_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G15gat), .B(G22gat), .Z(new_n311_));
  OAI21_X1  g110(.A(G1gat), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G15gat), .B(G22gat), .ZN(new_n313_));
  INV_X1    g112(.A(G1gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n305_), .A3(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n312_), .A2(new_n306_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n306_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n304_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n315_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G8gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n312_), .A2(new_n306_), .A3(new_n315_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n302_), .A2(new_n298_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G229gat), .A2(G233gat), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n318_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n322_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n324_), .B1(new_n327_), .B2(new_n323_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n286_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n323_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n324_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n318_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT76), .A3(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G113gat), .B(G141gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G169gat), .B(G197gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n329_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OR3_X1    g139(.A1(new_n325_), .A2(new_n328_), .A3(new_n337_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n329_), .A2(new_n334_), .A3(KEYINPUT77), .A4(new_n337_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n285_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n348_));
  AND2_X1   g147(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n349_));
  NOR2_X1   g148(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n348_), .B(G169gat), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT80), .B(G176gat), .ZN(new_n352_));
  INV_X1    g151(.A(G169gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT22), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n351_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(G169gat), .B1(new_n349_), .B2(new_n350_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT79), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n347_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(G183gat), .A3(G190gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G183gat), .ZN(new_n363_));
  INV_X1    g162(.A(G190gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT23), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371_));
  OR3_X1    g170(.A1(new_n347_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT25), .B(G183gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT26), .B(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n365_), .A2(new_n360_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n370_), .A2(new_n371_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n358_), .A2(new_n369_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT30), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G127gat), .B(G134gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G113gat), .B(G120gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n385_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G227gat), .A2(G233gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n389_), .B(KEYINPUT82), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT31), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n388_), .B(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G15gat), .B(G43gat), .Z(new_n393_));
  XOR2_X1   g192(.A(G71gat), .B(G99gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n392_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G197gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(G204gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT21), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT86), .B1(new_n397_), .B2(G204gat), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n400_), .B(new_n401_), .C1(new_n398_), .C2(new_n402_), .ZN(new_n403_));
  OR3_X1    g202(.A1(new_n397_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n404_));
  INV_X1    g203(.A(G204gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT85), .B1(new_n405_), .B2(G197gat), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n404_), .B(KEYINPUT21), .C1(new_n398_), .C2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G211gat), .B(G218gat), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n403_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT87), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n403_), .A2(new_n407_), .A3(KEYINPUT87), .A4(new_n409_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n402_), .A2(new_n398_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n397_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n408_), .B1(new_n417_), .B2(KEYINPUT88), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n400_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT21), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n418_), .A2(new_n421_), .A3(KEYINPUT89), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n401_), .B1(new_n417_), .B2(KEYINPUT88), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n409_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n414_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G155gat), .B(G162gat), .ZN(new_n428_));
  AND2_X1   g227(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G141gat), .A2(G148gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT2), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n430_), .B(KEYINPUT83), .ZN(new_n433_));
  AOI211_X1 g232(.A(new_n429_), .B(new_n432_), .C1(new_n433_), .C2(new_n431_), .ZN(new_n434_));
  INV_X1    g233(.A(G141gat), .ZN(new_n435_));
  INV_X1    g234(.A(G148gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n428_), .B1(new_n434_), .B2(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n428_), .A2(KEYINPUT1), .ZN(new_n441_));
  AND2_X1   g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n442_), .A2(KEYINPUT1), .B1(new_n435_), .B2(new_n436_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n433_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT29), .B1(new_n440_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n427_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G228gat), .A3(G233gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G228gat), .A2(G233gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n427_), .A2(new_n449_), .A3(new_n446_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G78gat), .B(G106gat), .Z(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT90), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n440_), .A2(KEYINPUT29), .A3(new_n445_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G22gat), .B(G50gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT28), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n454_), .B(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n448_), .A2(new_n450_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n451_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n452_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n458_), .A2(new_n462_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n385_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(new_n440_), .B2(new_n445_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n432_), .B1(new_n433_), .B2(new_n431_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n429_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n439_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n444_), .B(new_n385_), .C1(new_n470_), .C2(new_n428_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(KEYINPUT93), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT93), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n473_), .B(new_n466_), .C1(new_n440_), .C2(new_n445_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G225gat), .A2(G233gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n467_), .A2(KEYINPUT4), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(new_n474_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(KEYINPUT4), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n477_), .B1(new_n480_), .B2(new_n476_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G57gat), .B(G85gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(G1gat), .B(G29gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n481_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT33), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT33), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n481_), .A2(new_n490_), .A3(new_n487_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n381_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n427_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT89), .B1(new_n418_), .B2(new_n421_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n424_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n495_), .A2(new_n496_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n372_), .A2(new_n375_), .A3(KEYINPUT92), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n366_), .A2(new_n379_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n376_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT22), .B(G169gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n352_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n347_), .B1(new_n378_), .B2(new_n368_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n499_), .A2(new_n501_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n497_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G226gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT19), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AND4_X1   g308(.A1(KEYINPUT20), .A2(new_n494_), .A3(new_n506_), .A4(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT20), .B1(new_n427_), .B2(new_n493_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n497_), .A2(new_n381_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n497_), .A2(new_n505_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n513_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n510_), .B1(new_n517_), .B2(new_n508_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G8gat), .B(G36gat), .ZN(new_n519_));
  INV_X1    g318(.A(G92gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT18), .B(G64gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n518_), .A2(new_n524_), .ZN(new_n525_));
  AOI211_X1 g324(.A(new_n523_), .B(new_n510_), .C1(new_n517_), .C2(new_n508_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n480_), .A2(new_n476_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n528_), .B(new_n486_), .C1(new_n476_), .C2(new_n475_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n492_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n532_));
  OAI211_X1 g331(.A(G225gat), .B(G233gat), .C1(new_n532_), .C2(new_n478_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n486_), .A3(new_n477_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n524_), .A2(KEYINPUT32), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n488_), .A2(new_n534_), .B1(new_n518_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT91), .B1(new_n514_), .B2(KEYINPUT20), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT20), .ZN(new_n538_));
  AOI211_X1 g337(.A(new_n512_), .B(new_n538_), .C1(new_n497_), .C2(new_n381_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT95), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n540_), .A2(new_n541_), .A3(new_n509_), .A4(new_n516_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n513_), .A2(new_n515_), .A3(new_n509_), .A4(new_n516_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n494_), .A2(new_n506_), .A3(KEYINPUT20), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(new_n544_), .B2(new_n508_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n535_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT96), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n542_), .A2(new_n546_), .A3(KEYINPUT96), .A4(new_n547_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n536_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n465_), .B1(new_n530_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT27), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n523_), .B(KEYINPUT97), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n542_), .A2(new_n546_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n518_), .A2(new_n524_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(KEYINPUT27), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n488_), .A2(new_n534_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n561_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n396_), .B1(new_n553_), .B2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n560_), .A2(new_n465_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n396_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n561_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n345_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n320_), .A2(new_n321_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n571_), .A2(new_n218_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574_));
  INV_X1    g373(.A(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT16), .B(G183gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(new_n218_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n572_), .A2(new_n573_), .A3(new_n578_), .A4(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n572_), .A2(new_n579_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT74), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n578_), .A2(new_n573_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n580_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT75), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT75), .B(new_n580_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT68), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n264_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n248_), .A2(KEYINPUT68), .A3(new_n254_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n595_), .A2(new_n596_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n264_), .A2(new_n326_), .ZN(new_n598_));
  OAI211_X1 g397(.A(KEYINPUT35), .B(new_n593_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n304_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n602_));
  INV_X1    g401(.A(new_n598_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .A4(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n605_), .B(new_n606_), .Z(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(KEYINPUT36), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n599_), .A2(new_n604_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT71), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n599_), .A2(new_n604_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n607_), .B(KEYINPUT36), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT72), .Z(new_n616_));
  AND2_X1   g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n612_), .A2(new_n613_), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n613_), .B1(new_n612_), .B2(new_n618_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n590_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n568_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n561_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n314_), .A3(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n564_), .A2(new_n567_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n612_), .A2(new_n618_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n630_), .A2(new_n344_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n586_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n561_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n629_), .A2(new_n634_), .ZN(G1324gat));
  NAND3_X1  g434(.A1(new_n632_), .A2(new_n586_), .A3(new_n560_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n632_), .A2(KEYINPUT100), .A3(new_n586_), .A4(new_n560_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(G8gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n560_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n625_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n638_), .A2(new_n639_), .A3(G8gat), .A4(new_n641_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n643_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(G1325gat));
  OAI21_X1  g449(.A(G15gat), .B1(new_n633_), .B2(new_n396_), .ZN(new_n651_));
  XOR2_X1   g450(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n396_), .A2(G15gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n623_), .B2(new_n654_), .ZN(G1326gat));
  INV_X1    g454(.A(new_n465_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G22gat), .B1(new_n633_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT42), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(G22gat), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT104), .Z(new_n660_));
  OAI21_X1  g459(.A(new_n658_), .B1(new_n623_), .B2(new_n660_), .ZN(G1327gat));
  INV_X1    g460(.A(new_n590_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n619_), .A2(new_n620_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n536_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n509_), .B1(new_n540_), .B2(new_n516_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n523_), .B1(new_n665_), .B2(new_n510_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n558_), .A3(new_n529_), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT33), .B(new_n486_), .C1(new_n533_), .C2(new_n477_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n490_), .B1(new_n481_), .B2(new_n487_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n656_), .B1(new_n664_), .B2(new_n671_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n560_), .A2(new_n562_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n566_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NOR4_X1   g473(.A1(new_n396_), .A2(new_n560_), .A3(new_n465_), .A4(new_n626_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n663_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT43), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n663_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n680_), .A2(KEYINPUT105), .A3(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n344_), .B(new_n662_), .C1(new_n678_), .C2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n676_), .A2(new_n677_), .A3(KEYINPUT43), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n681_), .B1(new_n680_), .B2(KEYINPUT105), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n688_), .A2(KEYINPUT44), .A3(new_n344_), .A4(new_n662_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n685_), .A2(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(new_n626_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n590_), .A2(new_n631_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n568_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n626_), .A2(new_n287_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT106), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n691_), .A2(new_n287_), .B1(new_n693_), .B2(new_n695_), .ZN(G1328gat));
  NOR2_X1   g495(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n685_), .A2(new_n560_), .A3(new_n689_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G36gat), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n568_), .A2(new_n288_), .A3(new_n560_), .A4(new_n692_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n697_), .B1(new_n699_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n697_), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n705_), .B(new_n702_), .C1(new_n698_), .C2(G36gat), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1329gat));
  NAND4_X1  g506(.A1(new_n685_), .A2(G43gat), .A3(new_n566_), .A4(new_n689_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n294_), .B1(new_n693_), .B2(new_n396_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g510(.A1(new_n656_), .A2(new_n292_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n568_), .A2(new_n465_), .A3(new_n692_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n690_), .A2(new_n712_), .B1(new_n292_), .B2(new_n713_), .ZN(G1331gat));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n630_), .B2(new_n343_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n343_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT108), .B(new_n717_), .C1(new_n564_), .C2(new_n567_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n285_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n716_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n622_), .ZN(new_n721_));
  OR3_X1    g520(.A1(new_n721_), .A2(G57gat), .A3(new_n561_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n719_), .A2(new_n717_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n630_), .A2(new_n631_), .A3(new_n590_), .A4(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n561_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1332gat));
  OAI21_X1  g527(.A(G64gat), .B1(new_n724_), .B2(new_n644_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(KEYINPUT48), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT48), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n644_), .A2(G64gat), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n730_), .A2(new_n731_), .B1(new_n721_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT110), .ZN(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n724_), .B2(new_n396_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT49), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n396_), .A2(G71gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT111), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n721_), .B2(new_n738_), .ZN(G1334gat));
  OAI21_X1  g538(.A(G78gat), .B1(new_n724_), .B2(new_n656_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT50), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n656_), .A2(G78gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n721_), .B2(new_n742_), .ZN(G1335gat));
  AND2_X1   g542(.A1(new_n720_), .A2(new_n692_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G85gat), .B1(new_n744_), .B2(new_n626_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n285_), .A2(new_n343_), .A3(new_n662_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT112), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n626_), .A2(G85gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT113), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n745_), .B1(new_n748_), .B2(new_n750_), .ZN(G1336gat));
  AOI21_X1  g550(.A(G92gat), .B1(new_n744_), .B2(new_n560_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n748_), .A2(new_n560_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(G92gat), .B2(new_n753_), .ZN(G1337gat));
  NAND3_X1  g553(.A1(new_n744_), .A2(new_n566_), .A3(new_n237_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n748_), .A2(new_n566_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n756_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT114), .B1(new_n756_), .B2(G99gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n755_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT51), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n755_), .B(new_n761_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1338gat));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  AOI211_X1 g564(.A(new_n656_), .B(new_n747_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n764_), .B(new_n765_), .C1(new_n766_), .C2(new_n225_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n748_), .A2(new_n465_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n764_), .A2(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n768_), .A2(G106gat), .A3(new_n769_), .A4(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n720_), .A2(new_n225_), .A3(new_n465_), .A4(new_n692_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n767_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(G1339gat));
  NAND3_X1  g574(.A1(new_n565_), .A2(new_n566_), .A3(new_n626_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n586_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n631_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n248_), .A2(new_n217_), .A3(new_n254_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n271_), .B2(KEYINPUT12), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n217_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(KEYINPUT12), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n783_), .B2(new_n268_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n257_), .A2(new_n267_), .A3(new_n268_), .A4(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n785_), .A2(new_n786_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n257_), .A2(new_n267_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(KEYINPUT117), .A3(new_n270_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n257_), .A2(new_n267_), .A3(new_n268_), .A4(new_n789_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n784_), .A2(new_n791_), .A3(new_n793_), .A4(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n277_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(KEYINPUT56), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n343_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT119), .B1(new_n795_), .B2(new_n277_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n798_), .B(new_n799_), .C1(KEYINPUT56), .C2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n330_), .A2(new_n324_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n318_), .A2(new_n323_), .A3(new_n331_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n337_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n805_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n806_), .A2(new_n341_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n283_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n778_), .B1(new_n801_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT122), .B1(new_n810_), .B2(KEYINPUT57), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n799_), .B1(new_n800_), .B2(KEYINPUT56), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  AOI211_X1 g612(.A(KEYINPUT119), .B(new_n813_), .C1(new_n795_), .C2(new_n277_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n809_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  AND4_X1   g614(.A1(KEYINPUT122), .A2(new_n815_), .A3(KEYINPUT57), .A4(new_n631_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n811_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n796_), .A2(KEYINPUT56), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n795_), .A2(new_n813_), .A3(new_n277_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n818_), .A2(new_n281_), .A3(new_n808_), .A4(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT121), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT58), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(KEYINPUT121), .A3(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n663_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n815_), .A2(new_n631_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n777_), .B1(new_n817_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n621_), .A2(new_n285_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n343_), .ZN(new_n833_));
  NOR4_X1   g632(.A1(new_n621_), .A2(new_n285_), .A3(KEYINPUT54), .A4(new_n717_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n776_), .B1(new_n830_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837_), .B2(new_n717_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n828_), .B(new_n825_), .C1(new_n811_), .C2(new_n816_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n835_), .B1(new_n839_), .B2(new_n777_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT59), .B1(new_n840_), .B2(new_n776_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n776_), .A2(KEYINPUT59), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n820_), .A2(KEYINPUT121), .A3(new_n823_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n823_), .B1(new_n820_), .B2(KEYINPUT121), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n845_), .A2(new_n663_), .B1(new_n827_), .B2(new_n826_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n810_), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n590_), .B1(new_n846_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n842_), .B1(new_n851_), .B2(new_n835_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n841_), .A2(new_n717_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n838_), .B1(new_n853_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n719_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n837_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n841_), .A2(new_n285_), .A3(new_n852_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n855_), .ZN(G1341gat));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n586_), .B(new_n852_), .C1(new_n837_), .C2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G127gat), .ZN(new_n863_));
  NOR4_X1   g662(.A1(new_n840_), .A2(G127gat), .A3(new_n662_), .A4(new_n776_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n860_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  AOI211_X1 g665(.A(KEYINPUT123), .B(new_n864_), .C1(new_n862_), .C2(G127gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1342gat));
  AOI21_X1  g667(.A(G134gat), .B1(new_n837_), .B2(new_n778_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n841_), .A2(G134gat), .A3(new_n852_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n663_), .ZN(G1343gat));
  OR3_X1    g670(.A1(new_n840_), .A2(new_n656_), .A3(new_n566_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n644_), .A2(new_n626_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n872_), .A2(new_n343_), .A3(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n435_), .ZN(G1344gat));
  NOR3_X1   g674(.A1(new_n872_), .A2(new_n719_), .A3(new_n873_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT124), .B(G148gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1345gat));
  NOR3_X1   g677(.A1(new_n872_), .A2(new_n662_), .A3(new_n873_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n879_), .B(new_n881_), .ZN(G1346gat));
  NOR2_X1   g681(.A1(new_n872_), .A2(new_n873_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n883_), .A2(G162gat), .A3(new_n663_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G162gat), .B1(new_n883_), .B2(new_n778_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1347gat));
  NOR4_X1   g685(.A1(new_n644_), .A2(new_n396_), .A3(new_n626_), .A4(new_n465_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n851_), .B2(new_n835_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G169gat), .B1(new_n888_), .B2(new_n343_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n888_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n502_), .A3(new_n717_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n889_), .A2(new_n890_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n891_), .A2(new_n893_), .A3(new_n894_), .ZN(G1348gat));
  INV_X1    g694(.A(new_n887_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n840_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(G176gat), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n897_), .A2(new_n898_), .A3(new_n719_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n352_), .B1(new_n888_), .B2(new_n719_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n901_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n899_), .B1(new_n902_), .B2(new_n903_), .ZN(G1349gat));
  NOR3_X1   g703(.A1(new_n888_), .A2(new_n777_), .A3(new_n373_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n897_), .A2(new_n662_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n363_), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n888_), .B2(new_n679_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n778_), .A2(new_n374_), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n909_), .B(KEYINPUT126), .Z(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n888_), .B2(new_n910_), .ZN(G1351gat));
  NOR4_X1   g710(.A1(new_n840_), .A2(new_n562_), .A3(new_n644_), .A4(new_n566_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n717_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT127), .B1(new_n913_), .B2(new_n397_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n397_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n912_), .A2(new_n916_), .A3(G197gat), .A4(new_n717_), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n914_), .A2(new_n915_), .A3(new_n917_), .ZN(G1352gat));
  NAND2_X1  g717(.A1(new_n912_), .A2(new_n285_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n912_), .A2(new_n586_), .A3(new_n921_), .ZN(new_n922_));
  OR2_X1    g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1354gat));
  AOI21_X1  g723(.A(G218gat), .B1(new_n912_), .B2(new_n778_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n912_), .A2(G218gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n663_), .B2(new_n926_), .ZN(G1355gat));
endmodule


