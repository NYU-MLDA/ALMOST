//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G15gat), .B(G22gat), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  AND2_X1   g004(.A1(KEYINPUT71), .A2(G1gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT71), .A2(G1gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(G8gat), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n208_), .A2(KEYINPUT72), .A3(KEYINPUT14), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT72), .B1(new_n208_), .B2(KEYINPUT14), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n205_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n205_), .B(new_n212_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G29gat), .B(G36gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n217_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n214_), .A2(new_n215_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n203_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n208_), .A2(KEYINPUT14), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT72), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n208_), .A2(KEYINPUT72), .A3(KEYINPUT14), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n212_), .B1(new_n229_), .B2(new_n205_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n215_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n220_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n218_), .A2(KEYINPUT15), .A3(new_n219_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT15), .B1(new_n218_), .B2(new_n219_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(new_n215_), .A3(new_n214_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n236_), .A3(new_n202_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G113gat), .B(G141gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT75), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G169gat), .B(G197gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n224_), .A2(new_n237_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT76), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n224_), .A2(new_n237_), .A3(new_n245_), .A4(new_n242_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n224_), .A2(new_n237_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n241_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT77), .Z(new_n251_));
  INV_X1    g050(.A(KEYINPUT84), .ZN(new_n252_));
  NOR2_X1   g051(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G169gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT78), .B(KEYINPUT23), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(KEYINPUT80), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(G183gat), .A3(G190gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n262_), .A3(KEYINPUT23), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G183gat), .ZN(new_n265_));
  INV_X1    g064(.A(G190gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n255_), .B1(new_n268_), .B2(KEYINPUT81), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n259_), .A2(new_n263_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT81), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT25), .B(G183gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G190gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G169gat), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(KEYINPUT24), .A3(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n278_), .A2(KEYINPUT24), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n275_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n256_), .A2(new_n258_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT79), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT79), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n260_), .A2(new_n262_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(new_n286_), .A3(new_n289_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n269_), .A2(new_n272_), .B1(new_n282_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT30), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n282_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n272_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n254_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n292_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT83), .B1(new_n292_), .B2(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G227gat), .A2(G233gat), .ZN(new_n303_));
  INV_X1    g102(.A(G15gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G71gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT82), .B(G43gat), .ZN(new_n308_));
  INV_X1    g107(.A(G99gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n307_), .B(new_n310_), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n301_), .A2(new_n302_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(new_n311_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G127gat), .B(G134gat), .Z(new_n315_));
  XOR2_X1   g114(.A(G113gat), .B(G120gat), .Z(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT31), .Z(new_n318_));
  OR4_X1    g117(.A1(new_n252_), .A2(new_n312_), .A3(new_n314_), .A4(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n252_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n302_), .A2(new_n311_), .ZN(new_n321_));
  OAI211_X1 g120(.A(KEYINPUT84), .B(new_n313_), .C1(new_n321_), .C2(new_n301_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n322_), .A3(new_n318_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G197gat), .B(G204gat), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT21), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT21), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G211gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT87), .B1(new_n330_), .B2(G218gat), .ZN(new_n331_));
  INV_X1    g130(.A(G218gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(G211gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n326_), .A2(new_n329_), .A3(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n325_), .B(KEYINPUT21), .C1(new_n333_), .C2(new_n331_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n335_), .A2(KEYINPUT88), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT88), .B1(new_n335_), .B2(new_n336_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G228gat), .A2(G233gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT85), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n343_), .B1(new_n344_), .B2(KEYINPUT1), .ZN(new_n345_));
  OR2_X1    g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(KEYINPUT1), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n344_), .A2(new_n343_), .A3(KEYINPUT1), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n341_), .B(new_n342_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  OR3_X1    g149(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT2), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n342_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n350_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT86), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT86), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n350_), .A2(new_n360_), .A3(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n339_), .B(new_n340_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n335_), .A2(new_n336_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n358_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n365_), .B1(new_n366_), .B2(new_n363_), .ZN(new_n367_));
  AND2_X1   g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n371_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT89), .B1(new_n370_), .B2(new_n371_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n362_), .A2(new_n363_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G22gat), .B(G50gat), .Z(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT28), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n376_), .B(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n374_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n375_), .A2(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n373_), .A3(new_n372_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G85gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT0), .B(G57gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  NAND3_X1  g187(.A1(new_n359_), .A2(new_n361_), .A3(new_n317_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n317_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n366_), .A2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n389_), .A2(KEYINPUT4), .A3(new_n391_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT93), .B(KEYINPUT4), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n359_), .A2(new_n361_), .A3(new_n317_), .A4(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n388_), .B1(new_n395_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT94), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT94), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n404_), .A3(new_n401_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n255_), .B1(new_n290_), .B2(new_n267_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n282_), .A2(new_n264_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n365_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(KEYINPUT90), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n296_), .B2(new_n339_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n283_), .A2(KEYINPUT79), .B1(new_n287_), .B2(new_n288_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n415_), .A2(new_n286_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n411_), .B(new_n408_), .C1(new_n416_), .C2(new_n255_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT90), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n412_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT19), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(G8gat), .B(G36gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n365_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n431_), .A2(KEYINPUT20), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n365_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n335_), .A2(KEYINPUT88), .A3(new_n336_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n291_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(new_n422_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n424_), .A2(new_n430_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n430_), .B1(new_n424_), .B2(new_n438_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT92), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n424_), .A2(new_n438_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n429_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT92), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n439_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n400_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n396_), .A2(new_n393_), .A3(new_n398_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n388_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n447_), .A2(KEYINPUT33), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n406_), .A2(new_n442_), .A3(new_n446_), .A4(new_n450_), .ZN(new_n451_));
  OR3_X1    g250(.A1(new_n399_), .A2(new_n388_), .A3(new_n395_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n400_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n437_), .A2(KEYINPUT20), .A3(new_n423_), .A4(new_n431_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT95), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT95), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n432_), .A2(new_n456_), .A3(new_n423_), .A4(new_n437_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n414_), .A2(new_n417_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n422_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n455_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n429_), .A2(KEYINPUT32), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n443_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n453_), .B(new_n462_), .C1(new_n461_), .C2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n384_), .B1(new_n451_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n452_), .A2(new_n400_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(new_n382_), .A3(new_n380_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n460_), .A2(new_n430_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT96), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(new_n441_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n444_), .A2(KEYINPUT96), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT27), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT27), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n467_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n324_), .B1(new_n465_), .B2(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n319_), .A2(new_n466_), .A3(new_n323_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n472_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n477_), .B(new_n383_), .C1(new_n478_), .C2(new_n473_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n251_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G106gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n309_), .A2(new_n481_), .A3(KEYINPUT65), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT7), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT6), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(G99gat), .A3(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT7), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n489_), .A2(new_n309_), .A3(new_n481_), .A4(KEYINPUT65), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n483_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(G85gat), .A2(G92gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G85gat), .A2(G92gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT8), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G71gat), .B(G78gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT11), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n501_));
  INV_X1    g300(.A(new_n499_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n500_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n491_), .A2(KEYINPUT8), .A3(new_n494_), .ZN(new_n506_));
  XOR2_X1   g305(.A(KEYINPUT10), .B(G99gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT64), .B(G106gat), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n507_), .A2(new_n508_), .B1(new_n494_), .B2(KEYINPUT9), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT9), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n485_), .A2(new_n487_), .B1(new_n492_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n497_), .A2(new_n505_), .A3(new_n506_), .A4(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G230gat), .A2(G233gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT67), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT67), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n517_), .A3(new_n514_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n497_), .A2(new_n506_), .A3(new_n512_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n505_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n495_), .A2(new_n496_), .B1(new_n511_), .B2(new_n509_), .ZN(new_n523_));
  AOI211_X1 g322(.A(KEYINPUT12), .B(new_n505_), .C1(new_n523_), .C2(new_n506_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n516_), .B(new_n518_), .C1(new_n522_), .C2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n494_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT65), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n527_), .A2(G99gat), .A3(G106gat), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n528_), .A2(new_n489_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n526_), .B1(new_n529_), .B2(new_n483_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n512_), .B1(new_n530_), .B2(KEYINPUT8), .ZN(new_n531_));
  INV_X1    g330(.A(new_n506_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n521_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(KEYINPUT66), .A3(new_n513_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n514_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n520_), .A2(new_n536_), .A3(new_n521_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT5), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G176gat), .B(G204gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n525_), .A2(new_n538_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n525_), .B2(new_n538_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT68), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n518_), .B1(new_n524_), .B2(new_n522_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n516_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n538_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n542_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n525_), .A2(new_n538_), .A3(new_n543_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT68), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n554_));
  OR3_X1    g353(.A1(new_n547_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n554_), .B1(new_n547_), .B2(new_n553_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT36), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT34), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT35), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n520_), .B2(new_n221_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n520_), .A2(new_n235_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT69), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n566_), .A2(new_n567_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n570_), .B(new_n571_), .C1(new_n572_), .C2(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n572_), .B(new_n568_), .C1(new_n520_), .C2(new_n221_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n571_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n576_), .B(new_n573_), .C1(new_n577_), .C2(new_n569_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n563_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n578_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(KEYINPUT37), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n575_), .A2(new_n582_), .A3(new_n578_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n584_), .B(new_n586_), .C1(new_n581_), .C2(new_n563_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n230_), .A2(new_n231_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n505_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n591_), .B(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT73), .Z(new_n595_));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT16), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT74), .Z(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n594_), .A2(new_n603_), .A3(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n590_), .A2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n480_), .A2(new_n558_), .A3(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n466_), .A2(new_n207_), .A3(new_n206_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n583_), .B(KEYINPUT98), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n557_), .A2(new_n250_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(new_n605_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G1gat), .B1(new_n620_), .B2(new_n466_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n611_), .A2(new_n612_), .A3(new_n621_), .ZN(G1324gat));
  INV_X1    g421(.A(G8gat), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n478_), .A2(new_n473_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n607_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n619_), .A2(new_n624_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(G8gat), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(KEYINPUT39), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(KEYINPUT39), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n625_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g430(.A(new_n324_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n619_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G15gat), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n633_), .A2(KEYINPUT99), .A3(G15gat), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT41), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT41), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n640_), .A3(new_n637_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n607_), .A2(new_n304_), .A3(new_n632_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT100), .Z(new_n643_));
  NAND3_X1  g442(.A1(new_n639_), .A2(new_n641_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT101), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n639_), .A2(new_n646_), .A3(new_n643_), .A4(new_n641_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1326gat));
  INV_X1    g447(.A(G22gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n619_), .B2(new_n384_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT42), .Z(new_n651_));
  NAND3_X1  g450(.A1(new_n607_), .A2(new_n649_), .A3(new_n384_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1327gat));
  INV_X1    g452(.A(new_n605_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n617_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n476_), .A2(new_n479_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(new_n590_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n590_), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT43), .B(new_n659_), .C1(new_n476_), .C2(new_n479_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT44), .B(new_n655_), .C1(new_n658_), .C2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G29gat), .B1(new_n665_), .B2(new_n466_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n605_), .A2(new_n583_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT102), .Z(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n557_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n480_), .A2(new_n669_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n466_), .A2(G29gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n670_), .B2(new_n671_), .ZN(G1328gat));
  NOR4_X1   g471(.A1(new_n670_), .A2(G36gat), .A3(new_n473_), .A4(new_n478_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT45), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n663_), .A2(new_n624_), .A3(new_n664_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n663_), .A2(KEYINPUT103), .A3(new_n624_), .A4(new_n664_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G36gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n674_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n674_), .B(KEYINPUT46), .C1(new_n677_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1329gat));
  NAND4_X1  g483(.A1(new_n663_), .A2(G43gat), .A3(new_n632_), .A4(new_n664_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n670_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G43gat), .B1(new_n686_), .B2(new_n632_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(KEYINPUT104), .B2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n688_), .B1(KEYINPUT104), .B2(new_n685_), .ZN(new_n689_));
  XOR2_X1   g488(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n690_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n688_), .B(new_n692_), .C1(KEYINPUT104), .C2(new_n685_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1330gat));
  INV_X1    g493(.A(G50gat), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n665_), .A2(new_n695_), .A3(new_n383_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G50gat), .B1(new_n686_), .B2(new_n384_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1331gat));
  AND4_X1   g497(.A1(new_n251_), .A2(new_n615_), .A3(new_n557_), .A4(new_n654_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(G57gat), .A3(new_n453_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT108), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n657_), .A2(new_n250_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT106), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(new_n557_), .A3(new_n606_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n704_), .A2(KEYINPUT107), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(KEYINPUT107), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n453_), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n701_), .B1(new_n707_), .B2(new_n708_), .ZN(G1332gat));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n704_), .B(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(G64gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n624_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n699_), .B2(new_n624_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT48), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1333gat));
  NAND2_X1  g515(.A1(new_n632_), .A2(new_n306_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT109), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n711_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n306_), .B1(new_n699_), .B2(new_n632_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT49), .Z(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1334gat));
  INV_X1    g521(.A(G78gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n711_), .A2(new_n723_), .A3(new_n384_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n699_), .B2(new_n384_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT50), .Z(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1335gat));
  NOR2_X1   g526(.A1(new_n668_), .A2(new_n558_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n703_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G85gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n453_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n658_), .A2(new_n660_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n250_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n558_), .A2(new_n734_), .A3(new_n654_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n453_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n732_), .B1(new_n731_), .B2(new_n738_), .ZN(G1336gat));
  INV_X1    g538(.A(G92gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n730_), .A2(new_n740_), .A3(new_n624_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n624_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n740_), .B2(new_n743_), .ZN(G1337gat));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n632_), .A2(new_n507_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n729_), .B2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n309_), .B1(new_n736_), .B2(new_n632_), .ZN(new_n748_));
  OR3_X1    g547(.A1(new_n747_), .A2(new_n748_), .A3(KEYINPUT51), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT51), .B1(new_n747_), .B2(new_n748_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n733_), .A2(new_n384_), .A3(new_n735_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G106gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G106gat), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n384_), .A2(new_n508_), .ZN(new_n756_));
  OAI22_X1  g555(.A1(new_n754_), .A2(new_n755_), .B1(new_n729_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT53), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759_));
  OAI221_X1 g558(.A(new_n759_), .B1(new_n729_), .B2(new_n756_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1339gat));
  NAND3_X1  g560(.A1(new_n558_), .A2(new_n606_), .A3(new_n251_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n533_), .A2(KEYINPUT12), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n520_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n769_), .A2(KEYINPUT55), .A3(new_n516_), .A4(new_n518_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n513_), .B1(new_n524_), .B2(new_n522_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n535_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n766_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n542_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT111), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n773_), .A2(KEYINPUT111), .A3(new_n775_), .A4(new_n542_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n544_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n214_), .A2(new_n215_), .A3(new_n221_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n203_), .B1(new_n232_), .B2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n783_), .B2(new_n242_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n232_), .A2(new_n236_), .A3(new_n203_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n202_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT112), .A3(new_n241_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n786_), .A2(new_n788_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n547_), .B2(new_n553_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n780_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n583_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n784_), .A2(new_n788_), .A3(new_n785_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n247_), .A2(new_n552_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n774_), .A2(KEYINPUT56), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n773_), .A2(new_n775_), .A3(new_n542_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n798_), .A2(new_n799_), .A3(KEYINPUT58), .A4(new_n800_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n801_), .A2(new_n590_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n798_), .A2(new_n800_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n799_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n802_), .A2(new_n806_), .ZN(new_n807_));
  AND4_X1   g606(.A1(KEYINPUT113), .A2(new_n791_), .A3(KEYINPUT57), .A4(new_n792_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n583_), .B1(new_n780_), .B2(new_n790_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT113), .B1(new_n809_), .B2(KEYINPUT57), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n795_), .B(new_n807_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n654_), .B1(new_n811_), .B2(KEYINPUT114), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n806_), .A2(new_n802_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n813_), .B(new_n814_), .C1(new_n810_), .C2(new_n808_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n764_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n624_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(new_n453_), .A3(new_n383_), .A4(new_n632_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(G113gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n734_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n764_), .B1(new_n605_), .B2(new_n811_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT59), .B1(new_n818_), .B2(KEYINPUT115), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(KEYINPUT115), .B2(new_n818_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n819_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT116), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n825_), .B(new_n829_), .C1(new_n826_), .C2(new_n819_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n251_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n821_), .B1(new_n831_), .B2(new_n820_), .ZN(G1340gat));
  XNOR2_X1  g631(.A(KEYINPUT117), .B(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n827_), .B2(new_n558_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n557_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT118), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n819_), .B(new_n837_), .C1(new_n836_), .C2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n834_), .A2(new_n840_), .ZN(G1341gat));
  AOI21_X1  g640(.A(G127gat), .B1(new_n819_), .B2(new_n654_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n828_), .A2(new_n830_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n654_), .A2(G127gat), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT119), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n843_), .B2(new_n845_), .ZN(G1342gat));
  INV_X1    g645(.A(G134gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n819_), .A2(new_n847_), .A3(new_n614_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n659_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1343gat));
  NAND2_X1  g649(.A1(new_n384_), .A2(new_n453_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n624_), .A2(new_n632_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT120), .B1(new_n816_), .B2(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n762_), .B(KEYINPUT54), .ZN(new_n855_));
  INV_X1    g654(.A(new_n800_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n797_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT58), .B1(new_n857_), .B2(new_n799_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n801_), .A2(new_n590_), .ZN(new_n859_));
  OAI22_X1  g658(.A1(new_n858_), .A2(new_n859_), .B1(new_n809_), .B2(KEYINPUT57), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT113), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n809_), .A2(KEYINPUT113), .A3(KEYINPUT57), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n605_), .B1(new_n864_), .B2(new_n814_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n811_), .A2(KEYINPUT114), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n855_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n852_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n854_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n734_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n870_), .B2(new_n557_), .ZN(new_n874_));
  AOI211_X1 g673(.A(KEYINPUT122), .B(new_n558_), .C1(new_n854_), .C2(new_n869_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT121), .B(G148gat), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n874_), .A2(new_n875_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n868_), .B1(new_n867_), .B2(new_n852_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n811_), .A2(KEYINPUT114), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(new_n605_), .A3(new_n815_), .ZN(new_n881_));
  AOI211_X1 g680(.A(KEYINPUT120), .B(new_n853_), .C1(new_n881_), .C2(new_n855_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n557_), .B1(new_n879_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT122), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n870_), .A2(new_n873_), .A3(new_n557_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n876_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n878_), .A2(new_n886_), .ZN(G1345gat));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n870_), .B2(new_n654_), .ZN(new_n889_));
  AOI211_X1 g688(.A(KEYINPUT123), .B(new_n605_), .C1(new_n854_), .C2(new_n869_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n889_), .A2(new_n890_), .A3(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n654_), .B1(new_n879_), .B2(new_n882_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT123), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n870_), .A2(new_n888_), .A3(new_n654_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n891_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n893_), .A2(new_n897_), .ZN(G1346gat));
  AOI21_X1  g697(.A(G162gat), .B1(new_n870_), .B2(new_n614_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n590_), .A2(G162gat), .ZN(new_n900_));
  XOR2_X1   g699(.A(new_n900_), .B(KEYINPUT124), .Z(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n870_), .B2(new_n901_), .ZN(G1347gat));
  NAND2_X1  g701(.A1(new_n624_), .A2(new_n477_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n822_), .A2(new_n384_), .A3(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n734_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT62), .B1(new_n905_), .B2(KEYINPUT22), .ZN(new_n906_));
  OAI21_X1  g705(.A(G169gat), .B1(new_n905_), .B2(KEYINPUT62), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n276_), .B2(new_n906_), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n904_), .B2(new_n557_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n816_), .A2(new_n384_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n903_), .A2(new_n277_), .A3(new_n558_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(G1349gat));
  INV_X1    g712(.A(new_n904_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n914_), .A2(new_n273_), .A3(new_n605_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n911_), .A2(new_n624_), .A3(new_n477_), .A4(new_n654_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n265_), .B2(new_n916_), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n914_), .B2(new_n659_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n904_), .A2(new_n274_), .A3(new_n614_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1351gat));
  NAND3_X1  g719(.A1(new_n324_), .A2(new_n466_), .A3(new_n384_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n624_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n816_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n734_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n557_), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT126), .B(G204gat), .Z(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1353gat));
  NAND2_X1  g729(.A1(new_n925_), .A2(new_n654_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT63), .B(G211gat), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n931_), .A2(new_n934_), .A3(new_n330_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n931_), .A2(KEYINPUT127), .A3(new_n934_), .A4(new_n330_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n933_), .B1(new_n937_), .B2(new_n938_), .ZN(G1354gat));
  NAND3_X1  g738(.A1(new_n925_), .A2(new_n332_), .A3(new_n614_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n925_), .A2(new_n590_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(new_n332_), .ZN(G1355gat));
endmodule


