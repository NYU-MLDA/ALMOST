//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n210_), .A2(KEYINPUT81), .A3(KEYINPUT22), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT22), .B1(new_n210_), .B2(KEYINPUT81), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n204_), .A2(new_n206_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n210_), .A2(new_n212_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(KEYINPUT24), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n218_), .A2(new_n219_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n215_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n224_), .B(KEYINPUT30), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT82), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(KEYINPUT82), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G15gat), .B(G43gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G71gat), .B(G99gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  MUX2_X1   g031(.A(new_n226_), .B(new_n227_), .S(new_n232_), .Z(new_n233_));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234_));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT31), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n233_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT85), .ZN(new_n239_));
  OR2_X1    g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G155gat), .A2(G162gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(G141gat), .B2(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(G141gat), .ZN(new_n245_));
  INV_X1    g044(.A(G148gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(KEYINPUT3), .ZN(new_n247_));
  AND3_X1   g046(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT84), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n244_), .A2(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G141gat), .A2(G148gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n251_), .A2(KEYINPUT84), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n242_), .B1(new_n250_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n245_), .A2(new_n246_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n256_), .A2(new_n252_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n240_), .A2(new_n259_), .A3(new_n241_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n239_), .B1(new_n255_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n247_), .A2(new_n244_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n248_), .A2(new_n249_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n254_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n242_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n258_), .A2(new_n260_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(KEYINPUT85), .A3(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n262_), .A2(new_n269_), .A3(new_n236_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n265_), .A2(new_n266_), .B1(new_n260_), .B2(new_n258_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n234_), .B(new_n235_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT97), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n262_), .A2(new_n269_), .A3(KEYINPUT97), .A4(new_n236_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT4), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n270_), .A2(KEYINPUT4), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G1gat), .B(G29gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT0), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(G57gat), .Z(new_n286_));
  INV_X1    g085(.A(G85gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n281_), .A2(new_n282_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n238_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G226gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT19), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT20), .ZN(new_n298_));
  INV_X1    g097(.A(G211gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(G218gat), .ZN(new_n300_));
  INV_X1    g099(.A(G218gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(G211gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT87), .B1(new_n300_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(G211gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(G218gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT87), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(G197gat), .A2(G204gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G197gat), .A2(G204gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(KEYINPUT21), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT21), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n308_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n306_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT88), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n303_), .A2(new_n320_), .A3(new_n307_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n311_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT89), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT89), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n319_), .A2(new_n321_), .A3(new_n325_), .A4(new_n322_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n316_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT93), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n217_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n217_), .A2(new_n328_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n216_), .A3(new_n330_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT22), .B(G169gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n212_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n331_), .A2(new_n332_), .B1(new_n209_), .B2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n298_), .B1(new_n327_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n311_), .B1(new_n308_), .B2(KEYINPUT88), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n325_), .B1(new_n337_), .B2(new_n321_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n326_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n315_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT94), .B1(new_n340_), .B2(new_n224_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT94), .ZN(new_n342_));
  INV_X1    g141(.A(new_n224_), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n327_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n297_), .B(new_n336_), .C1(new_n341_), .C2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT20), .B1(new_n327_), .B2(new_n335_), .ZN(new_n346_));
  AOI211_X1 g145(.A(new_n316_), .B(new_n224_), .C1(new_n324_), .C2(new_n326_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n296_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G64gat), .B(G92gat), .Z(new_n350_));
  XNOR2_X1  g149(.A(G8gat), .B(G36gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n349_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT96), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n345_), .A2(new_n354_), .A3(new_n348_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT27), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n345_), .A2(KEYINPUT96), .A3(new_n354_), .A4(new_n348_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n262_), .A2(new_n269_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n363_), .A2(KEYINPUT29), .ZN(new_n364_));
  XOR2_X1   g163(.A(G22gat), .B(G50gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT28), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n364_), .B(new_n366_), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT92), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n367_), .A2(KEYINPUT92), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT86), .Z(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n327_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n363_), .A2(KEYINPUT29), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT90), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT90), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n377_), .A3(new_n374_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n255_), .B2(new_n261_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n372_), .B1(new_n327_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n379_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n381_), .B1(new_n379_), .B2(new_n385_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n368_), .B(new_n369_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n388_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n390_), .A2(KEYINPUT92), .A3(new_n367_), .A4(new_n386_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT101), .ZN(new_n393_));
  INV_X1    g192(.A(new_n346_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n347_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n297_), .A3(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n315_), .B(new_n335_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT20), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n342_), .B1(new_n327_), .B2(new_n343_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n340_), .A2(KEYINPUT94), .A3(new_n224_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n396_), .B1(new_n401_), .B2(new_n297_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n393_), .B1(new_n402_), .B2(new_n355_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n358_), .A2(KEYINPUT27), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n393_), .A3(new_n355_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT102), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n358_), .A2(KEYINPUT27), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n346_), .A2(new_n296_), .A3(new_n347_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n336_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(new_n296_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT101), .B1(new_n411_), .B2(new_n354_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n408_), .A2(new_n412_), .A3(KEYINPUT102), .A4(new_n406_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n362_), .B(new_n392_), .C1(new_n407_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT103), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n408_), .A2(new_n412_), .A3(new_n406_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT102), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n345_), .A2(new_n354_), .A3(new_n348_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n354_), .B1(new_n345_), .B2(new_n348_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n421_), .A2(new_n422_), .A3(KEYINPUT96), .ZN(new_n423_));
  INV_X1    g222(.A(new_n361_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n420_), .A2(new_n413_), .B1(new_n425_), .B2(new_n360_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(KEYINPUT103), .A3(new_n392_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n294_), .B1(new_n417_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n238_), .B(KEYINPUT83), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n281_), .A2(new_n282_), .A3(new_n290_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n290_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n354_), .A2(KEYINPUT32), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n345_), .A2(new_n348_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n411_), .B2(new_n433_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT100), .B1(new_n432_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT100), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n402_), .A2(KEYINPUT32), .A3(new_n354_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n292_), .A2(new_n437_), .A3(new_n438_), .A4(new_n434_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT98), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n291_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n281_), .A2(KEYINPUT98), .A3(new_n282_), .A4(new_n290_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT99), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n359_), .A2(new_n361_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n442_), .A2(KEYINPUT99), .A3(new_n443_), .A4(new_n444_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n277_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n290_), .B1(new_n279_), .B2(new_n276_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n430_), .A2(KEYINPUT33), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .A4(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n440_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n392_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n420_), .A2(new_n413_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n389_), .A2(new_n391_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n362_), .A4(new_n432_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n429_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n428_), .A2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G29gat), .B(G36gat), .Z(new_n461_));
  XOR2_X1   g260(.A(G43gat), .B(G50gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT15), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465_));
  INV_X1    g264(.A(G1gat), .ZN(new_n466_));
  INV_X1    g265(.A(G8gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT14), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n464_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n463_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n473_), .A2(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n472_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n473_), .B(new_n471_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n479_), .A2(KEYINPUT79), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(KEYINPUT79), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n476_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G169gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G197gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT80), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n482_), .B(new_n486_), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n460_), .A2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G57gat), .B(G64gat), .Z(new_n490_));
  INV_X1    g289(.A(KEYINPUT11), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n491_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT68), .B(G71gat), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G78gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT68), .B(G71gat), .ZN(new_n497_));
  INV_X1    g296(.A(G78gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n494_), .A2(new_n496_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT69), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n500_), .A2(KEYINPUT69), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n493_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n500_), .A2(KEYINPUT69), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(new_n492_), .A3(new_n501_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(new_n471_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G231gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G127gat), .B(G155gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G183gat), .B(G211gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT17), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n517_), .A2(KEYINPUT77), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519_));
  OR3_X1    g318(.A1(new_n510_), .A2(new_n519_), .A3(new_n515_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(KEYINPUT77), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n522_), .B(KEYINPUT78), .Z(new_n523_));
  INV_X1    g322(.A(KEYINPUT74), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G190gat), .B(G218gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G134gat), .B(G162gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n527_), .B(KEYINPUT36), .Z(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT73), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT34), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT9), .ZN(new_n534_));
  INV_X1    g333(.A(G92gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n287_), .B2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G85gat), .B(G92gat), .Z(new_n537_));
  OAI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(new_n534_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT65), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT6), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(G106gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT10), .B(G99gat), .Z(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT8), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n540_), .B(KEYINPUT6), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT66), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT66), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n542_), .A2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT7), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n537_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n547_), .B1(new_n555_), .B2(KEYINPUT67), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n557_), .A3(new_n537_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n537_), .A2(new_n547_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n548_), .B2(new_n553_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n463_), .B(new_n546_), .C1(new_n559_), .C2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n546_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n545_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n538_), .A2(KEYINPUT65), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n538_), .A2(KEYINPUT65), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT70), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n561_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n464_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  AOI211_X1 g371(.A(new_n530_), .B(new_n533_), .C1(new_n562_), .C2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n532_), .A2(KEYINPUT35), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n533_), .A2(new_n530_), .ZN(new_n575_));
  AND4_X1   g374(.A1(new_n574_), .A2(new_n562_), .A3(new_n572_), .A4(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n529_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n562_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(KEYINPUT35), .A3(new_n532_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n527_), .A2(KEYINPUT36), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n562_), .A2(new_n572_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n524_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n577_), .B2(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT74), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n528_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n585_), .A2(KEYINPUT75), .A3(new_n587_), .A4(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT75), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n586_), .B2(KEYINPUT74), .ZN(new_n592_));
  AOI211_X1 g391(.A(new_n524_), .B(new_n584_), .C1(new_n577_), .C2(new_n582_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n570_), .A2(new_n571_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n507_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n502_), .A2(new_n493_), .A3(new_n503_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n492_), .B1(new_n505_), .B2(new_n501_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n571_), .B2(new_n568_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n596_), .A2(new_n598_), .B1(new_n602_), .B2(new_n597_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT64), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n571_), .A2(new_n568_), .ZN(new_n607_));
  AOI211_X1 g406(.A(KEYINPUT71), .B(new_n606_), .C1(new_n607_), .C2(new_n507_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT71), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n546_), .B(new_n507_), .C1(new_n559_), .C2(new_n561_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n610_), .B2(new_n605_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n603_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n602_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n606_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(G120gat), .B(G148gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT72), .B(G204gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT5), .B(G176gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n615_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n620_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(new_n614_), .A3(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(KEYINPUT13), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(KEYINPUT13), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n523_), .A2(new_n595_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n489_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n489_), .A2(KEYINPUT104), .A3(new_n628_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n631_), .A2(new_n466_), .A3(new_n292_), .A4(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n588_), .A2(new_n582_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n460_), .A2(new_n523_), .A3(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n627_), .A2(new_n488_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n432_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n633_), .A2(new_n634_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n641_), .A3(new_n642_), .ZN(G1324gat));
  OAI21_X1  g442(.A(G8gat), .B1(new_n640_), .B2(new_n426_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT105), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n426_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n631_), .A2(new_n467_), .A3(new_n648_), .A4(new_n632_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n644_), .A2(new_n645_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT105), .B(G8gat), .C1(new_n640_), .C2(new_n426_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(KEYINPUT39), .A3(new_n653_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n650_), .A2(new_n651_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n651_), .B1(new_n650_), .B2(new_n654_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1325gat));
  INV_X1    g456(.A(new_n429_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G15gat), .B1(new_n640_), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT41), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n631_), .A2(new_n632_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n661_), .A2(G15gat), .A3(new_n658_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n640_), .B2(new_n392_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n392_), .A2(G22gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n661_), .B2(new_n666_), .ZN(G1327gat));
  XNOR2_X1  g466(.A(new_n522_), .B(KEYINPUT78), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n668_), .A2(new_n627_), .A3(new_n636_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n489_), .A2(new_n669_), .ZN(new_n670_));
  OR3_X1    g469(.A1(new_n670_), .A2(G29gat), .A3(new_n432_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n415_), .A2(new_n416_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT103), .B1(new_n426_), .B2(new_n392_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n293_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n458_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n457_), .B1(new_n440_), .B2(new_n453_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n658_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n672_), .B1(new_n679_), .B2(new_n595_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n672_), .B(new_n595_), .C1(new_n428_), .C2(new_n459_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n523_), .B(new_n639_), .C1(new_n680_), .C2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT107), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n590_), .A2(new_n594_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT43), .B1(new_n460_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n681_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n523_), .A4(new_n639_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n684_), .A2(new_n685_), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n639_), .ZN(new_n692_));
  AOI211_X1 g491(.A(new_n668_), .B(new_n692_), .C1(new_n687_), .C2(new_n681_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n432_), .B1(new_n693_), .B2(KEYINPUT44), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(new_n694_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n695_), .A2(KEYINPUT108), .A3(G29gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT108), .B1(new_n695_), .B2(G29gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n671_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  INV_X1    g497(.A(new_n670_), .ZN(new_n699_));
  INV_X1    g498(.A(G36gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n648_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT45), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n426_), .B1(new_n693_), .B2(KEYINPUT44), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n691_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT46), .B(new_n702_), .C1(new_n704_), .C2(new_n700_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n701_), .B(KEYINPUT45), .Z(new_n707_));
  AOI21_X1  g506(.A(new_n700_), .B1(new_n691_), .B2(new_n703_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(G1329gat));
  INV_X1    g509(.A(G43gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n238_), .B1(new_n693_), .B2(KEYINPUT44), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n691_), .B2(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n670_), .A2(G43gat), .A3(new_n658_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT47), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  INV_X1    g515(.A(new_n714_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n688_), .A2(KEYINPUT44), .A3(new_n523_), .A4(new_n639_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n238_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n683_), .B2(KEYINPUT107), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n690_), .B2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n716_), .B(new_n717_), .C1(new_n722_), .C2(new_n711_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n715_), .A2(new_n723_), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n699_), .B2(new_n457_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n718_), .A2(G50gat), .A3(new_n457_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n691_), .ZN(G1331gat));
  NAND2_X1  g526(.A1(new_n627_), .A2(new_n488_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n638_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(G57gat), .A3(new_n292_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n732_), .A2(new_n733_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n460_), .A2(new_n728_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n523_), .A2(new_n595_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G57gat), .B1(new_n739_), .B2(new_n292_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n734_), .A2(new_n735_), .A3(new_n740_), .ZN(G1332gat));
  INV_X1    g540(.A(G64gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n742_), .A3(new_n648_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n731_), .B2(new_n648_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n745_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(KEYINPUT48), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT48), .B1(new_n746_), .B2(new_n747_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n743_), .B1(new_n748_), .B2(new_n749_), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n730_), .B2(new_n658_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT49), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n658_), .A2(G71gat), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT111), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n738_), .B2(new_n754_), .ZN(G1334gat));
  OAI21_X1  g554(.A(G78gat), .B1(new_n730_), .B2(new_n392_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n739_), .A2(new_n498_), .A3(new_n457_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT112), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n757_), .A2(new_n761_), .A3(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n668_), .A2(new_n636_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n736_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT113), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n736_), .A2(new_n767_), .A3(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n287_), .A3(new_n292_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n688_), .A2(KEYINPUT114), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n688_), .A2(KEYINPUT114), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n728_), .A2(new_n668_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(new_n292_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n770_), .B1(new_n775_), .B2(new_n287_), .ZN(G1336gat));
  AOI21_X1  g575(.A(G92gat), .B1(new_n769_), .B2(new_n648_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n777_), .A2(KEYINPUT115), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(KEYINPUT115), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n648_), .A2(G92gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT116), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n778_), .A2(new_n779_), .B1(new_n774_), .B2(new_n781_), .ZN(G1337gat));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(KEYINPUT118), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n771_), .A2(new_n429_), .A3(new_n772_), .A4(new_n773_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(G99gat), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n719_), .A2(new_n544_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT117), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n784_), .B1(new_n787_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n790_), .B(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n786_), .C1(KEYINPUT118), .C2(new_n783_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n795_), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n769_), .A2(new_n543_), .A3(new_n457_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n688_), .A2(new_n457_), .A3(new_n523_), .A4(new_n729_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n612_), .A2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n603_), .B(KEYINPUT55), .C1(new_n608_), .C2(new_n611_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n603_), .A2(new_n610_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n606_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n806_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n620_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT56), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n812_), .A3(new_n620_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n811_), .A2(new_n487_), .A3(new_n623_), .A4(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n624_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n472_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n477_), .A2(new_n475_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n485_), .A3(new_n817_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT120), .Z(new_n819_));
  OR2_X1    g618(.A1(new_n482_), .A2(new_n485_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT121), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n815_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n637_), .B1(new_n814_), .B2(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT57), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n811_), .A2(new_n623_), .A3(new_n822_), .A4(new_n813_), .ZN(new_n826_));
  XOR2_X1   g625(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n595_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT123), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n826_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n830_), .B1(new_n826_), .B2(new_n831_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n829_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n523_), .B1(new_n825_), .B2(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n625_), .A2(new_n626_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n487_), .B1(KEYINPUT119), .B2(KEYINPUT54), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n837_), .A2(new_n668_), .A3(new_n686_), .A4(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n839_), .B(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n836_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n238_), .B1(new_n417_), .B2(new_n427_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n292_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT59), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n432_), .B1(new_n836_), .B2(new_n843_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n845_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n488_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n488_), .A2(G113gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n846_), .B2(new_n853_), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT60), .B1(new_n627_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n627_), .B1(new_n846_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(G120gat), .B1(new_n851_), .B2(new_n857_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n846_), .A2(new_n856_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(KEYINPUT60), .B2(new_n859_), .ZN(G1341gat));
  OAI21_X1  g659(.A(G127gat), .B1(new_n851_), .B2(new_n523_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n523_), .A2(G127gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n846_), .B2(new_n862_), .ZN(G1342gat));
  OAI21_X1  g662(.A(G134gat), .B1(new_n851_), .B2(new_n686_), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n636_), .A2(G134gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n846_), .B2(new_n865_), .ZN(G1343gat));
  NAND4_X1  g665(.A1(new_n848_), .A2(new_n426_), .A3(new_n457_), .A4(new_n658_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n488_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n245_), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n837_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n246_), .ZN(G1345gat));
  NOR2_X1   g670(.A1(new_n867_), .A2(new_n523_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n872_), .B(new_n874_), .ZN(G1346gat));
  OAI21_X1  g674(.A(G162gat), .B1(new_n867_), .B2(new_n686_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n636_), .A2(G162gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n867_), .B2(new_n877_), .ZN(G1347gat));
  NOR3_X1   g677(.A1(new_n658_), .A2(new_n426_), .A3(new_n292_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n844_), .A2(new_n392_), .A3(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G169gat), .B1(new_n880_), .B2(new_n488_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n880_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(new_n487_), .A3(new_n333_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n881_), .A2(new_n882_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n885_), .A3(new_n886_), .ZN(G1348gat));
  NOR2_X1   g686(.A1(new_n837_), .A2(new_n212_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(new_n844_), .B2(new_n392_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n824_), .A2(KEYINPUT57), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n892_), .B(new_n637_), .C1(new_n814_), .C2(new_n823_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n686_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n834_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n832_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n668_), .B1(new_n894_), .B2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n839_), .B(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n889_), .B(new_n392_), .C1(new_n898_), .C2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n879_), .B(new_n888_), .C1(new_n890_), .C2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT125), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n392_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT124), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n901_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n879_), .A4(new_n888_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n212_), .B1(new_n880_), .B2(new_n837_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n904_), .A2(new_n909_), .A3(new_n910_), .ZN(G1349gat));
  NOR3_X1   g710(.A1(new_n880_), .A2(new_n216_), .A3(new_n523_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n907_), .A2(new_n668_), .A3(new_n879_), .ZN(new_n913_));
  INV_X1    g712(.A(G183gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n880_), .B2(new_n686_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n637_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n880_), .B2(new_n917_), .ZN(G1351gat));
  NAND3_X1  g717(.A1(new_n658_), .A2(new_n457_), .A3(new_n432_), .ZN(new_n919_));
  AOI211_X1 g718(.A(new_n426_), .B(new_n919_), .C1(new_n836_), .C2(new_n843_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n487_), .ZN(new_n921_));
  INV_X1    g720(.A(G197gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT126), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n922_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n921_), .A2(KEYINPUT126), .A3(new_n922_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1352gat));
  NAND2_X1  g726(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT127), .B(G204gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n920_), .A2(new_n627_), .ZN(new_n930_));
  MUX2_X1   g729(.A(new_n928_), .B(new_n929_), .S(new_n930_), .Z(G1353gat));
  NAND2_X1  g730(.A1(new_n920_), .A2(new_n668_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  AND2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n932_), .B2(new_n933_), .ZN(G1354gat));
  NAND3_X1  g735(.A1(new_n920_), .A2(new_n301_), .A3(new_n637_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n920_), .A2(new_n595_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n937_), .B1(new_n939_), .B2(new_n301_), .ZN(G1355gat));
endmodule


