//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT80), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n202_), .B(new_n203_), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n205_), .B1(new_n206_), .B2(KEYINPUT80), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G71gat), .B(G99gat), .ZN(new_n208_));
  INV_X1    g007(.A(G43gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT30), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT25), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G183gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT76), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT26), .B(G190gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT75), .B(G183gat), .Z(new_n217_));
  OAI211_X1 g016(.A(new_n215_), .B(new_n216_), .C1(new_n213_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT77), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n218_), .A2(new_n225_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT78), .B(G169gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n220_), .B1(G190gat), .B2(new_n217_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n229_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G227gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT79), .B(G15gat), .Z(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n237_), .A2(new_n238_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n212_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n235_), .B(new_n236_), .Z(new_n243_));
  INV_X1    g042(.A(new_n238_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(new_n211_), .A3(new_n239_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(KEYINPUT81), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT31), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT31), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n242_), .A2(KEYINPUT81), .A3(new_n249_), .A4(new_n246_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n207_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n248_), .A2(new_n207_), .A3(new_n250_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G106gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G141gat), .ZN(new_n258_));
  INV_X1    g057(.A(G148gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G155gat), .ZN(new_n262_));
  INV_X1    g061(.A(G162gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n262_), .A2(new_n263_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT82), .ZN(new_n268_));
  INV_X1    g067(.A(new_n265_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(KEYINPUT1), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n257_), .B(new_n261_), .C1(new_n268_), .C2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT83), .B1(new_n261_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n260_), .A2(new_n274_), .A3(KEYINPUT2), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n273_), .B(new_n275_), .C1(new_n260_), .C2(KEYINPUT2), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n256_), .B(KEYINPUT3), .Z(new_n277_));
  OAI211_X1 g076(.A(new_n269_), .B(new_n264_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n271_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT29), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G197gat), .A2(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT86), .B(G197gat), .ZN(new_n282_));
  OAI211_X1 g081(.A(KEYINPUT21), .B(new_n281_), .C1(new_n282_), .C2(G204gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(G211gat), .B(G218gat), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G204gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G197gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n283_), .B(new_n285_), .C1(new_n288_), .C2(KEYINPUT21), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT21), .A3(new_n284_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n280_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G228gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT85), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n294_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n291_), .B(KEYINPUT87), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n280_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n295_), .A2(G78gat), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(G78gat), .B1(new_n295_), .B2(new_n298_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n255_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n295_), .A2(new_n298_), .ZN(new_n302_));
  INV_X1    g101(.A(G78gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n295_), .A2(G78gat), .A3(new_n298_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(G106gat), .A3(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n306_), .A3(KEYINPUT84), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G22gat), .B(G50gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n279_), .A2(KEYINPUT29), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n308_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n301_), .A2(new_n306_), .A3(KEYINPUT84), .A4(new_n313_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n309_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n254_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n309_), .A2(new_n314_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n312_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n309_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n248_), .A2(new_n207_), .A3(new_n250_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n322_), .A2(new_n251_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n317_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n216_), .B(KEYINPUT89), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT25), .B(G183gat), .Z(new_n327_));
  OAI211_X1 g126(.A(new_n225_), .B(new_n227_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n220_), .B1(G183gat), .B2(G190gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT22), .B(G169gat), .Z(new_n330_));
  OAI211_X1 g129(.A(new_n329_), .B(new_n226_), .C1(G176gat), .C2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n291_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n333_), .B(KEYINPUT20), .C1(new_n291_), .C2(new_n235_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT19), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n332_), .A2(new_n291_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT20), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n235_), .B2(new_n291_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT18), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G64gat), .ZN(new_n345_));
  INV_X1    g144(.A(G92gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n338_), .A2(new_n342_), .A3(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n350_), .A2(KEYINPUT27), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n334_), .A2(new_n336_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n341_), .B1(new_n297_), .B2(new_n332_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n352_), .B1(new_n336_), .B2(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(KEYINPUT94), .B(new_n349_), .C1(new_n354_), .C2(new_n347_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n349_), .A2(KEYINPUT94), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n351_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n279_), .A2(new_n207_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n271_), .A2(new_n278_), .A3(new_n206_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT4), .B1(new_n279_), .B2(new_n207_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n362_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n365_), .B2(KEYINPUT4), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n363_), .B1(new_n366_), .B2(new_n361_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(G85gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT0), .ZN(new_n370_));
  INV_X1    g169(.A(G57gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n372_), .B(new_n363_), .C1(new_n366_), .C2(new_n361_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n359_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n325_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT90), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n348_), .A2(new_n379_), .A3(new_n349_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n367_), .A2(new_n373_), .ZN(new_n383_));
  MUX2_X1   g182(.A(new_n365_), .B(new_n366_), .S(new_n361_), .Z(new_n384_));
  AOI22_X1  g183(.A1(new_n383_), .A2(KEYINPUT33), .B1(new_n384_), .B2(new_n373_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT91), .B(KEYINPUT33), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n375_), .A2(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n387_), .A2(KEYINPUT92), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(KEYINPUT92), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n382_), .B(new_n385_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n338_), .A2(new_n342_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(KEYINPUT93), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(KEYINPUT32), .B2(new_n347_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT93), .B1(new_n338_), .B2(new_n342_), .ZN(new_n394_));
  AND4_X1   g193(.A1(KEYINPUT32), .A2(new_n354_), .A3(new_n347_), .A4(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n376_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  AND4_X1   g196(.A1(new_n321_), .A2(new_n397_), .A3(new_n320_), .A4(new_n254_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n378_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT12), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT11), .ZN(new_n402_));
  AND2_X1   g201(.A1(G57gat), .A2(G64gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G57gat), .A2(G64gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT66), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G64gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n371_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT66), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G57gat), .A2(G64gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n402_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G71gat), .B(G78gat), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n411_), .B(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n405_), .A2(new_n410_), .A3(new_n402_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n401_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT67), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT7), .ZN(new_n418_));
  INV_X1    g217(.A(G99gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n255_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G99gat), .A2(G106gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n346_), .A2(G85gat), .ZN(new_n427_));
  INV_X1    g226(.A(G85gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(G92gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT8), .B1(new_n426_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT10), .B(G99gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n423_), .A2(new_n425_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT9), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n433_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n438_), .A2(new_n435_), .A3(G92gat), .A4(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n431_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n424_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT65), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n434_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT65), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n420_), .A2(new_n446_), .A3(new_n424_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n430_), .A2(KEYINPUT8), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n417_), .B1(new_n441_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n431_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n432_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n255_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n436_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n445_), .A4(new_n440_), .ZN(new_n456_));
  AND4_X1   g255(.A1(new_n417_), .A2(new_n450_), .A3(new_n452_), .A4(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n416_), .B1(new_n451_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n456_), .A3(new_n452_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n403_), .A2(new_n404_), .A3(KEYINPUT66), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n408_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT11), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n413_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n411_), .A2(new_n412_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n415_), .A3(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT12), .B1(new_n459_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n459_), .A2(new_n465_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G230gat), .A2(G233gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n458_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n467_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n459_), .A2(new_n465_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G120gat), .B(G148gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT5), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(G176gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G204gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n470_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT68), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT68), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n470_), .A2(new_n481_), .A3(new_n474_), .A4(new_n478_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n478_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n470_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n474_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n484_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT69), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n489_), .A2(KEYINPUT13), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(KEYINPUT13), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n488_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n490_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(G29gat), .A2(G36gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G29gat), .A2(G36gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n209_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n209_), .A3(new_n497_), .ZN(new_n500_));
  AOI21_X1  g299(.A(G50gat), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n500_), .ZN(new_n502_));
  INV_X1    g301(.A(G50gat), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n498_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT15), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  INV_X1    g309(.A(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G8gat), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n515_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n509_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n505_), .A2(new_n517_), .A3(new_n516_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n501_), .A2(new_n504_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n518_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n521_), .B1(new_n524_), .B2(new_n520_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G113gat), .B(G141gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n221_), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n529_), .B(G197gat), .Z(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(KEYINPUT73), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n530_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n523_), .A2(new_n518_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(new_n509_), .B2(new_n518_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n525_), .B1(new_n534_), .B2(new_n521_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT73), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n532_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT74), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n495_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G232gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT34), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT70), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n459_), .A2(new_n523_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n459_), .A2(KEYINPUT67), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n441_), .A2(new_n417_), .A3(new_n450_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI211_X1 g349(.A(new_n546_), .B(new_n547_), .C1(new_n550_), .C2(new_n509_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n543_), .A2(new_n544_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n545_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(KEYINPUT35), .A3(new_n542_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(G134gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(new_n263_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n558_), .A2(new_n559_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n554_), .B(new_n555_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n555_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n560_), .B1(new_n564_), .B2(new_n553_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT37), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT16), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G183gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(G211gat), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n465_), .B(new_n518_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT71), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n576_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT72), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n579_), .B2(new_n576_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n583_), .B(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n571_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n400_), .A2(KEYINPUT95), .A3(new_n540_), .A4(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n377_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n317_), .B2(new_n324_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n540_), .B(new_n587_), .C1(new_n590_), .C2(new_n398_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n511_), .A3(new_n376_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT38), .ZN(new_n596_));
  INV_X1    g395(.A(new_n495_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n538_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n586_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n566_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n590_), .B2(new_n398_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT96), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n605_), .B(new_n602_), .C1(new_n590_), .C2(new_n398_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n601_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(new_n376_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n596_), .B1(new_n511_), .B2(new_n608_), .ZN(G1324gat));
  NAND4_X1  g408(.A1(new_n588_), .A2(new_n593_), .A3(new_n512_), .A4(new_n359_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT97), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n613_));
  INV_X1    g412(.A(new_n359_), .ZN(new_n614_));
  AOI211_X1 g413(.A(new_n614_), .B(new_n601_), .C1(new_n604_), .C2(new_n606_), .ZN(new_n615_));
  OAI211_X1 g414(.A(KEYINPUT98), .B(new_n613_), .C1(new_n615_), .C2(new_n512_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n607_), .A2(new_n359_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n613_), .A2(KEYINPUT98), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(KEYINPUT98), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n617_), .A2(G8gat), .A3(new_n618_), .A4(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n612_), .A2(new_n616_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n612_), .A2(new_n622_), .A3(new_n616_), .A4(new_n620_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1325gat));
  INV_X1    g425(.A(KEYINPUT41), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n607_), .A2(new_n323_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(G15gat), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n629_), .B1(new_n628_), .B2(G15gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n627_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(KEYINPUT41), .A3(new_n630_), .ZN(new_n635_));
  INV_X1    g434(.A(G15gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n594_), .A2(new_n636_), .A3(new_n323_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n637_), .A2(new_n638_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n633_), .A2(new_n635_), .A3(new_n639_), .A4(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n315_), .A2(new_n316_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n594_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n607_), .A2(new_n644_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(G22gat), .ZN(new_n648_));
  AOI211_X1 g447(.A(KEYINPUT42), .B(new_n642_), .C1(new_n607_), .C2(new_n644_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(G1327gat));
  NAND3_X1  g449(.A1(new_n400_), .A2(new_n566_), .A3(new_n586_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n540_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n376_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n571_), .B1(new_n590_), .B2(new_n398_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT43), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n657_), .B(new_n571_), .C1(new_n590_), .C2(new_n398_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n659_), .A2(KEYINPUT44), .A3(new_n599_), .A4(new_n586_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(G29gat), .A3(new_n376_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n659_), .A2(new_n599_), .A3(new_n586_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n654_), .B1(new_n661_), .B2(new_n664_), .ZN(G1328gat));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n359_), .A3(new_n660_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G36gat), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n359_), .B(KEYINPUT102), .Z(new_n669_));
  NAND3_X1  g468(.A1(new_n653_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n653_), .A2(new_n668_), .A3(new_n673_), .A4(new_n669_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n667_), .A2(KEYINPUT46), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n614_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n668_), .B1(new_n678_), .B2(new_n660_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n672_), .A2(new_n674_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n676_), .A2(new_n681_), .ZN(G1329gat));
  NAND2_X1  g481(.A1(new_n653_), .A2(new_n323_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n209_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n664_), .A2(new_n323_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n660_), .A2(G43gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT105), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n684_), .B(new_n689_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1330gat));
  AOI21_X1  g492(.A(G50gat), .B1(new_n653_), .B2(new_n644_), .ZN(new_n694_));
  AOI211_X1 g493(.A(new_n503_), .B(new_n643_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n660_), .ZN(G1331gat));
  NAND2_X1  g495(.A1(new_n587_), .A2(new_n495_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT106), .ZN(new_n698_));
  INV_X1    g497(.A(new_n538_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n400_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n376_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n371_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT107), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n604_), .A2(new_n606_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n600_), .A2(new_n539_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n495_), .A3(new_n705_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n706_), .A2(new_n371_), .A3(new_n701_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n703_), .A2(new_n707_), .ZN(G1332gat));
  INV_X1    g507(.A(new_n700_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(new_n406_), .A3(new_n669_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n669_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n706_), .A2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT109), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n712_), .A2(G64gat), .A3(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n712_), .B2(G64gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n710_), .B1(new_n715_), .B2(new_n716_), .ZN(G1333gat));
  OR3_X1    g516(.A1(new_n700_), .A2(G71gat), .A3(new_n254_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n704_), .A2(new_n323_), .A3(new_n495_), .A4(new_n705_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G71gat), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT111), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(new_n722_), .A3(G71gat), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n721_), .A2(new_n723_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n718_), .B1(new_n726_), .B2(new_n727_), .ZN(G1334gat));
  NAND3_X1  g527(.A1(new_n709_), .A2(new_n303_), .A3(new_n644_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n704_), .A2(new_n644_), .A3(new_n495_), .A4(new_n705_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(G78gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n730_), .B2(G78gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT112), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(new_n729_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1335gat));
  NOR2_X1   g537(.A1(new_n597_), .A2(new_n538_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n651_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n376_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT113), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n659_), .A2(new_n586_), .A3(new_n739_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n376_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n743_), .B1(new_n745_), .B2(new_n746_), .ZN(G1336gat));
  AOI21_X1  g546(.A(G92gat), .B1(new_n741_), .B2(new_n359_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n711_), .A2(new_n346_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n745_), .B2(new_n749_), .ZN(G1337gat));
  OAI21_X1  g549(.A(G99gat), .B1(new_n744_), .B2(new_n254_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n741_), .A2(new_n453_), .A3(new_n323_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  OR2_X1    g553(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(G1338gat));
  NAND3_X1  g555(.A1(new_n741_), .A2(new_n255_), .A3(new_n644_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n659_), .A2(new_n644_), .A3(new_n586_), .A4(new_n739_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G106gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT53), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n757_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1339gat));
  INV_X1    g565(.A(G113gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n469_), .B1(new_n458_), .B2(new_n468_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT116), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n550_), .A2(new_n416_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n771_), .B(KEYINPUT55), .C1(new_n772_), .C2(new_n469_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n770_), .A2(new_n470_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n470_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n484_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT56), .B(new_n484_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n534_), .A2(new_n521_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n524_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n532_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n535_), .B2(new_n532_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n483_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT58), .B1(new_n780_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n788_), .B(new_n785_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n787_), .A2(new_n789_), .A3(new_n570_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n483_), .A2(new_n538_), .A3(KEYINPUT115), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT115), .B1(new_n483_), .B2(new_n538_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n466_), .A2(new_n467_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n465_), .A2(KEYINPUT12), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n471_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n771_), .B1(new_n797_), .B2(KEYINPUT55), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n768_), .A2(KEYINPUT116), .A3(new_n769_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n485_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n770_), .A2(new_n470_), .A3(new_n773_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n484_), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n777_), .B(new_n478_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n793_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n488_), .A2(new_n784_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT57), .B1(new_n807_), .B2(new_n602_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n790_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(KEYINPUT57), .A3(new_n602_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n600_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n600_), .A2(new_n597_), .A3(new_n539_), .A4(new_n570_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n324_), .A2(new_n701_), .A3(new_n359_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n767_), .B1(new_n818_), .B2(new_n699_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n819_), .A2(KEYINPUT117), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(KEYINPUT117), .ZN(new_n821_));
  INV_X1    g620(.A(new_n817_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT59), .B1(new_n815_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n767_), .A2(KEYINPUT120), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n767_), .A2(KEYINPUT120), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n539_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT119), .B1(new_n790_), .B2(new_n808_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n780_), .A2(new_n793_), .B1(new_n488_), .B2(new_n784_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n566_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n786_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n788_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n780_), .A2(KEYINPUT58), .A3(new_n786_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n571_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n830_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n827_), .A2(new_n810_), .A3(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n814_), .B1(new_n837_), .B2(new_n586_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n817_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n823_), .B(new_n826_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n820_), .A2(new_n821_), .A3(new_n841_), .ZN(G1340gat));
  INV_X1    g641(.A(new_n818_), .ZN(new_n843_));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n597_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n843_), .B(new_n845_), .C1(KEYINPUT60), .C2(new_n844_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n823_), .B(new_n495_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n848_), .B2(new_n844_), .ZN(G1341gat));
  INV_X1    g648(.A(G127gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n814_), .A2(new_n600_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n822_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT121), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n586_), .A2(new_n850_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n823_), .B(new_n854_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1342gat));
  INV_X1    g655(.A(G134gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n818_), .B2(new_n602_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n570_), .A2(new_n857_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n823_), .B(new_n859_), .C1(new_n840_), .C2(new_n838_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT122), .ZN(G1343gat));
  NOR3_X1   g661(.A1(new_n815_), .A2(new_n701_), .A3(new_n317_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n711_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n699_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n258_), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n597_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(new_n259_), .ZN(G1345gat));
  NOR2_X1   g667(.A1(new_n864_), .A2(new_n586_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT61), .B(G155gat), .Z(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  NOR3_X1   g670(.A1(new_n864_), .A2(new_n263_), .A3(new_n570_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n864_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n566_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n263_), .B2(new_n874_), .ZN(G1347gat));
  NOR3_X1   g674(.A1(new_n711_), .A2(new_n376_), .A3(new_n324_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT123), .B1(new_n838_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  INV_X1    g678(.A(new_n810_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n830_), .A2(new_n834_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(KEYINPUT119), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n600_), .B1(new_n882_), .B2(new_n836_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n879_), .B(new_n876_), .C1(new_n883_), .C2(new_n814_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n699_), .A2(new_n330_), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(KEYINPUT124), .Z(new_n886_));
  NAND3_X1  g685(.A1(new_n878_), .A2(new_n884_), .A3(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n538_), .B(new_n876_), .C1(new_n883_), .C2(new_n814_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n888_), .A2(new_n889_), .A3(G169gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n888_), .B2(G169gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n887_), .B1(new_n890_), .B2(new_n891_), .ZN(G1348gat));
  NAND3_X1  g691(.A1(new_n878_), .A2(new_n495_), .A3(new_n884_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n222_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n816_), .A2(G176gat), .A3(new_n495_), .A4(new_n876_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n894_), .A2(KEYINPUT125), .A3(new_n895_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1349gat));
  NAND4_X1  g699(.A1(new_n878_), .A2(new_n327_), .A3(new_n884_), .A4(new_n600_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n217_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n877_), .B2(new_n851_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n878_), .A2(new_n571_), .A3(new_n884_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G190gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n602_), .A2(new_n326_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n878_), .A2(new_n884_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1351gat));
  NOR2_X1   g708(.A1(new_n815_), .A2(new_n317_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n711_), .A2(new_n376_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n699_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT126), .B(G197gat), .Z(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1352gat));
  NOR2_X1   g714(.A1(new_n912_), .A2(new_n597_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(KEYINPUT127), .B2(new_n286_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT127), .B(G204gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n916_), .B2(new_n918_), .ZN(G1353gat));
  NOR2_X1   g718(.A1(new_n912_), .A2(new_n586_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  AND2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n923_), .B1(new_n920_), .B2(new_n921_), .ZN(G1354gat));
  INV_X1    g723(.A(new_n912_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n925_), .A2(G218gat), .A3(new_n571_), .ZN(new_n926_));
  AOI21_X1  g725(.A(G218gat), .B1(new_n925_), .B2(new_n566_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1355gat));
endmodule


