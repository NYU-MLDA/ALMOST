//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n597_, new_n598_, new_n599_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT69), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT69), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(new_n204_), .A3(new_n206_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT74), .B(G1gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n214_), .A2(G8gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT14), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n213_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G1gat), .B(G8gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n210_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n219_), .B(new_n221_), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n220_), .A2(new_n225_), .B1(new_n226_), .B2(new_n224_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G113gat), .B(G141gat), .Z(new_n228_));
  XNOR2_X1  g027(.A(G169gat), .B(G197gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n230_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G127gat), .B(G134gat), .Z(new_n235_));
  XOR2_X1   g034(.A(G113gat), .B(G120gat), .Z(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT31), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(G15gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT22), .ZN(new_n244_));
  OAI21_X1  g043(.A(G169gat), .B1(new_n244_), .B2(KEYINPUT80), .ZN(new_n245_));
  INV_X1    g044(.A(G176gat), .ZN(new_n246_));
  INV_X1    g045(.A(G169gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT22), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n245_), .B(new_n246_), .C1(KEYINPUT80), .C2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT81), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(KEYINPUT81), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G183gat), .A2(G190gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT23), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(G183gat), .B2(G190gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(new_n253_), .A3(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT78), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT24), .A3(new_n250_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT79), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n259_), .A2(new_n262_), .A3(KEYINPUT24), .A4(new_n250_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n259_), .A2(KEYINPUT24), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT25), .B(G183gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G190gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n267_), .A2(new_n255_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n261_), .A2(new_n263_), .A3(new_n264_), .A4(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G71gat), .B(G99gat), .ZN(new_n270_));
  INV_X1    g069(.A(G43gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n257_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n257_), .B2(new_n269_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n243_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n276_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(new_n242_), .A3(new_n274_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n239_), .B1(new_n280_), .B2(KEYINPUT82), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT83), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT82), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n277_), .A2(new_n279_), .A3(new_n283_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n281_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT83), .B1(new_n280_), .B2(new_n238_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n284_), .B2(new_n281_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G64gat), .B(G92gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT92), .ZN(new_n290_));
  XOR2_X1   g089(.A(G8gat), .B(G36gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G226gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT19), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT22), .B(G169gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n246_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n256_), .A2(new_n250_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT89), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n256_), .A2(new_n301_), .A3(new_n250_), .A4(new_n298_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n258_), .A2(new_n303_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n260_), .A2(new_n255_), .A3(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n266_), .B(KEYINPUT88), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n265_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n300_), .A2(new_n302_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G197gat), .A2(G204gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT86), .B(G204gat), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n309_), .B1(new_n310_), .B2(G197gat), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n311_), .A2(KEYINPUT21), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G211gat), .B(G218gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n310_), .A2(G197gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT21), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(G197gat), .B2(G204gat), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n314_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n313_), .A2(new_n316_), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n312_), .A2(new_n318_), .B1(new_n311_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT20), .B1(new_n308_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n257_), .A2(new_n320_), .A3(new_n269_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n296_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT90), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT20), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n300_), .A2(new_n302_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n305_), .A2(new_n307_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n320_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n326_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n322_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT90), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(new_n296_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n325_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n296_), .ZN(new_n336_));
  OAI211_X1 g135(.A(KEYINPUT20), .B(new_n336_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n320_), .B1(new_n257_), .B2(new_n269_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n294_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n294_), .ZN(new_n342_));
  AOI211_X1 g141(.A(new_n342_), .B(new_n339_), .C1(new_n325_), .C2(new_n334_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT1), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(G155gat), .A3(G162gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT85), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n355_), .B1(new_n356_), .B2(KEYINPUT1), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(KEYINPUT84), .B2(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n357_), .A2(KEYINPUT84), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n351_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n349_), .B(KEYINPUT3), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n347_), .B(KEYINPUT2), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n356_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n355_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n360_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n237_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n237_), .B1(new_n360_), .B2(new_n366_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(KEYINPUT4), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n358_), .A2(new_n359_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n350_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n368_), .B1(new_n373_), .B2(new_n365_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT93), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT93), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n370_), .A2(new_n377_), .A3(KEYINPUT4), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n346_), .B(new_n371_), .C1(new_n376_), .C2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n369_), .A2(new_n370_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n345_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G1gat), .B(G29gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G57gat), .B(G85gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n384_), .B(new_n385_), .Z(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n379_), .A2(new_n381_), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT33), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n380_), .B2(new_n346_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n371_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(new_n346_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n344_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n294_), .A2(KEYINPUT32), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n328_), .A2(new_n320_), .A3(new_n299_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT20), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n296_), .B1(new_n396_), .B2(new_n338_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n331_), .A2(new_n336_), .A3(new_n322_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n394_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n339_), .B1(new_n325_), .B2(new_n334_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(new_n394_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n379_), .A2(new_n381_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n386_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n388_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n330_), .B1(new_n367_), .B2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(G228gat), .A3(G233gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n410_), .B(new_n330_), .C1(new_n367_), .C2(new_n407_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n406_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n409_), .A2(new_n411_), .A3(new_n406_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n367_), .A2(new_n407_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G22gat), .B(G50gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT28), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n416_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT87), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n419_), .B1(new_n412_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n415_), .A2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n413_), .A2(new_n420_), .A3(new_n414_), .A4(new_n419_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n401_), .A2(new_n404_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n288_), .B1(new_n393_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n404_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n400_), .A2(new_n294_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n398_), .A2(new_n397_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n426_), .B1(new_n430_), .B2(new_n342_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n427_), .A2(new_n428_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n422_), .A2(new_n423_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n425_), .A2(new_n436_), .A3(KEYINPUT95), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n427_), .A2(new_n432_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n438_), .A2(new_n434_), .A3(new_n428_), .A4(new_n288_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n425_), .A2(new_n436_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT95), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n234_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G230gat), .A2(G233gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G57gat), .B(G64gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G71gat), .B(G78gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT11), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(KEYINPUT11), .ZN(new_n450_));
  INV_X1    g249(.A(new_n448_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n447_), .A2(KEYINPUT11), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G92gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(KEYINPUT9), .ZN(new_n456_));
  AND2_X1   g255(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G99gat), .A2(G106gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT6), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(G99gat), .A3(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n465_));
  INV_X1    g264(.A(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G85gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n455_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G85gat), .A2(G92gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(KEYINPUT9), .A3(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n459_), .A2(new_n464_), .A3(new_n468_), .A4(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT65), .ZN(new_n474_));
  INV_X1    g273(.A(G99gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n466_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT7), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n474_), .A2(new_n478_), .A3(new_n475_), .A4(new_n466_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n464_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n470_), .A2(new_n471_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n454_), .B(new_n473_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT66), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n482_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT8), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT66), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n454_), .A4(new_n473_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n473_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(new_n454_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n446_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT12), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n495_), .B2(new_n454_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n446_), .B1(new_n495_), .B2(new_n454_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT12), .B(new_n449_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n483_), .A2(new_n484_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n464_), .A2(new_n472_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n504_), .A2(KEYINPUT67), .A3(new_n468_), .A4(new_n459_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT67), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n473_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n502_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n499_), .A2(new_n500_), .A3(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n497_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G120gat), .B(G148gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT5), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G176gat), .B(G204gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n511_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n517_), .B1(new_n521_), .B2(KEYINPUT13), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G231gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n454_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(new_n219_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G127gat), .B(G155gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT76), .ZN(new_n528_));
  XOR2_X1   g327(.A(G183gat), .B(G211gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n526_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT77), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n526_), .A2(new_n534_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(KEYINPUT17), .A2(new_n533_), .B1(new_n535_), .B2(new_n532_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n535_), .A2(KEYINPUT17), .A3(new_n532_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n505_), .A2(new_n507_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n490_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n212_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n495_), .A2(new_n210_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(new_n544_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n543_), .B(new_n548_), .C1(new_n544_), .C2(new_n547_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT36), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT71), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n556_), .A2(KEYINPUT36), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n551_), .A2(new_n552_), .A3(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n540_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT72), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n561_), .B1(new_n559_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT72), .B1(new_n553_), .B2(new_n558_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT37), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n540_), .B(KEYINPUT37), .C1(new_n566_), .C2(new_n567_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n444_), .A2(new_n523_), .A3(new_n539_), .A4(new_n572_), .ZN(new_n573_));
  OR3_X1    g372(.A1(new_n573_), .A2(new_n428_), .A3(new_n214_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n575_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n562_), .B(KEYINPUT97), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n523_), .A2(new_n233_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(new_n538_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G1gat), .B1(new_n582_), .B2(new_n428_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n576_), .A2(new_n577_), .A3(new_n583_), .ZN(G1324gat));
  OR3_X1    g383(.A1(new_n573_), .A2(G8gat), .A3(new_n438_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G8gat), .B1(new_n582_), .B2(new_n438_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n586_), .A2(KEYINPUT39), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(KEYINPUT39), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n585_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT40), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(G1325gat));
  INV_X1    g390(.A(new_n288_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G15gat), .B1(new_n582_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT41), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n573_), .A2(G15gat), .A3(new_n592_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(G1326gat));
  OAI21_X1  g395(.A(G22gat), .B1(new_n582_), .B2(new_n434_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT42), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n434_), .A2(G22gat), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n598_), .B1(new_n573_), .B2(new_n599_), .ZN(G1327gat));
  NAND2_X1  g399(.A1(new_n578_), .A2(new_n538_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n523_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n444_), .A2(KEYINPUT101), .A3(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n443_), .A2(new_n439_), .A3(new_n437_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(new_n233_), .A3(new_n603_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n604_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n428_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(G29gat), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n580_), .A2(new_n539_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n569_), .A2(new_n614_), .A3(new_n570_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n613_), .B1(new_n605_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n571_), .A2(new_n613_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n620_));
  OAI211_X1 g419(.A(KEYINPUT44), .B(new_n612_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT100), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n437_), .A2(new_n439_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT95), .B1(new_n425_), .B2(new_n436_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n617_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT43), .ZN(new_n626_));
  INV_X1    g425(.A(new_n619_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n605_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(KEYINPUT44), .A4(new_n612_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n622_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n612_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT99), .B(KEYINPUT44), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n404_), .A2(G29gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n611_), .B1(new_n637_), .B2(new_n638_), .ZN(G1328gat));
  INV_X1    g438(.A(KEYINPUT46), .ZN(new_n640_));
  INV_X1    g439(.A(G36gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n438_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n632_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n438_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n604_), .A2(new_n608_), .A3(new_n641_), .A4(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT45), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n640_), .B1(new_n643_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n645_), .B(KEYINPUT45), .ZN(new_n649_));
  INV_X1    g448(.A(new_n612_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n644_), .B1(new_n651_), .B2(new_n634_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n622_), .B2(new_n631_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n649_), .B(KEYINPUT46), .C1(new_n653_), .C2(new_n641_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n648_), .A2(new_n654_), .ZN(G1329gat));
  NOR2_X1   g454(.A1(new_n592_), .A2(new_n271_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n630_), .B1(new_n651_), .B2(KEYINPUT44), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n625_), .A2(KEYINPUT43), .B1(new_n605_), .B2(new_n627_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  NOR4_X1   g458(.A1(new_n658_), .A2(KEYINPUT100), .A3(new_n659_), .A4(new_n650_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n636_), .B(new_n656_), .C1(new_n657_), .C2(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(KEYINPUT102), .B(G43gat), .Z(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n609_), .B2(new_n592_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT47), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(new_n666_), .A3(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1330gat));
  INV_X1    g467(.A(G50gat), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n434_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n636_), .B(new_n670_), .C1(new_n657_), .C2(new_n660_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n669_), .B1(new_n609_), .B2(new_n434_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT103), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n675_), .A3(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1331gat));
  NAND2_X1  g476(.A1(new_n605_), .A2(new_n234_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT104), .Z(new_n679_));
  NOR3_X1   g478(.A1(new_n571_), .A2(new_n523_), .A3(new_n538_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n404_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682_));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n681_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n682_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n523_), .A2(new_n233_), .A3(new_n538_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n579_), .A2(new_n686_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n687_), .A2(new_n683_), .A3(new_n428_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT106), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n684_), .A2(new_n685_), .A3(new_n689_), .ZN(G1332gat));
  OAI21_X1  g489(.A(G64gat), .B1(new_n687_), .B2(new_n438_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT48), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n679_), .A2(new_n680_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n438_), .A2(G64gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(new_n693_), .B2(new_n694_), .ZN(G1333gat));
  OAI21_X1  g494(.A(G71gat), .B1(new_n687_), .B2(new_n592_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT49), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n592_), .A2(G71gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n693_), .B2(new_n698_), .ZN(G1334gat));
  OAI21_X1  g498(.A(G78gat), .B1(new_n687_), .B2(new_n434_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(KEYINPUT108), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(KEYINPUT108), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n704_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n701_), .A2(new_n702_), .A3(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n434_), .A2(G78gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT109), .ZN(new_n709_));
  OAI22_X1  g508(.A1(new_n705_), .A2(new_n707_), .B1(new_n693_), .B2(new_n709_), .ZN(G1335gat));
  NOR3_X1   g509(.A1(new_n523_), .A2(new_n233_), .A3(new_n539_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n629_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n404_), .B1(new_n458_), .B2(new_n457_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n601_), .A2(new_n523_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n679_), .A2(new_n404_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n469_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT110), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(new_n719_), .A3(new_n469_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n714_), .B1(new_n718_), .B2(new_n720_), .ZN(G1336gat));
  OAI21_X1  g520(.A(G92gat), .B1(new_n712_), .B2(new_n438_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n679_), .A2(new_n715_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n644_), .A2(new_n455_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT111), .ZN(G1337gat));
  OAI21_X1  g525(.A(G99gat), .B1(new_n712_), .B2(new_n592_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n288_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n723_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g529(.A1(new_n679_), .A2(new_n466_), .A3(new_n435_), .A4(new_n715_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n629_), .A2(new_n435_), .A3(new_n711_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(G106gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G106gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n731_), .B(new_n737_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1339gat));
  INV_X1    g540(.A(KEYINPUT59), .ZN(new_n742_));
  NOR4_X1   g541(.A1(new_n644_), .A2(new_n435_), .A3(new_n428_), .A4(new_n592_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT120), .Z(new_n744_));
  NAND2_X1  g543(.A1(new_n511_), .A2(new_n516_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n220_), .B(new_n224_), .C1(new_n219_), .C2(new_n221_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n230_), .B1(new_n226_), .B2(new_n223_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(new_n232_), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT114), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n473_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n454_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT12), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n501_), .B1(new_n541_), .B2(new_n490_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n485_), .A2(new_n445_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n754_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n750_), .A2(KEYINPUT114), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n751_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n510_), .A2(KEYINPUT114), .A3(new_n750_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n499_), .A2(new_n486_), .A3(new_n492_), .A4(new_n509_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n761_), .A2(KEYINPUT115), .A3(new_n446_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT115), .B1(new_n761_), .B2(new_n446_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n759_), .B(new_n760_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT116), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n761_), .A2(new_n446_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n761_), .A2(KEYINPUT115), .A3(new_n446_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n510_), .A2(KEYINPUT114), .A3(new_n750_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n751_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n758_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n510_), .B2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n771_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n770_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n765_), .A2(new_n777_), .A3(new_n515_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n765_), .A2(new_n777_), .A3(KEYINPUT56), .A4(new_n515_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n749_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n571_), .B1(KEYINPUT58), .B2(new_n782_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n782_), .A2(KEYINPUT58), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n517_), .A2(new_n232_), .A3(new_n748_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n781_), .A2(KEYINPUT117), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n516_), .B1(new_n764_), .B2(KEYINPUT116), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(KEYINPUT56), .A4(new_n777_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n780_), .A3(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n233_), .A2(new_n745_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n786_), .B1(new_n793_), .B2(KEYINPUT118), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n795_), .A3(new_n792_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n578_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n785_), .B1(new_n797_), .B2(KEYINPUT57), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n791_), .A2(new_n795_), .A3(new_n792_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n795_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n786_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n799_), .B1(new_n802_), .B2(new_n578_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n539_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n538_), .A2(new_n233_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT113), .Z(new_n806_));
  NOR3_X1   g605(.A1(new_n806_), .A2(new_n602_), .A3(new_n571_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT54), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n742_), .B(new_n744_), .C1(new_n804_), .C2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n744_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT119), .B1(new_n797_), .B2(KEYINPUT57), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n812_), .B(new_n799_), .C1(new_n802_), .C2(new_n578_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n798_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n538_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n808_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n810_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n233_), .B(new_n809_), .C1(new_n817_), .C2(new_n742_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G113gat), .ZN(new_n819_));
  INV_X1    g618(.A(G113gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n820_), .A3(new_n233_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1340gat));
  OAI211_X1 g621(.A(new_n602_), .B(new_n809_), .C1(new_n817_), .C2(new_n742_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT121), .B(G120gat), .Z(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n523_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n817_), .B(new_n827_), .C1(KEYINPUT60), .C2(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1341gat));
  NAND2_X1  g628(.A1(new_n817_), .A2(new_n539_), .ZN(new_n830_));
  INV_X1    g629(.A(G127gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n539_), .B2(KEYINPUT122), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(KEYINPUT122), .B2(new_n831_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n809_), .B(new_n834_), .C1(new_n817_), .C2(new_n742_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n832_), .A2(new_n835_), .ZN(G1342gat));
  OAI211_X1 g635(.A(new_n571_), .B(new_n809_), .C1(new_n817_), .C2(new_n742_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G134gat), .ZN(new_n838_));
  INV_X1    g637(.A(G134gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n817_), .A2(new_n839_), .A3(new_n578_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1343gat));
  NAND2_X1  g640(.A1(new_n815_), .A2(new_n816_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n288_), .A2(new_n434_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n644_), .A2(new_n428_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n842_), .A2(new_n233_), .A3(new_n843_), .A4(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g645(.A1(new_n842_), .A2(new_n602_), .A3(new_n843_), .A4(new_n844_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT123), .B(G148gat), .Z(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1345gat));
  NAND4_X1  g648(.A1(new_n842_), .A2(new_n539_), .A3(new_n843_), .A4(new_n844_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT61), .B(G155gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1346gat));
  INV_X1    g651(.A(new_n843_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n854_), .A2(new_n844_), .ZN(new_n855_));
  INV_X1    g654(.A(G162gat), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n615_), .A2(new_n616_), .A3(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n578_), .A3(new_n844_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n855_), .A2(new_n857_), .B1(new_n858_), .B2(new_n856_), .ZN(G1347gat));
  NOR2_X1   g658(.A1(new_n438_), .A2(new_n404_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n288_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n435_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n233_), .B(new_n862_), .C1(new_n804_), .C2(new_n808_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n863_), .A2(KEYINPUT125), .A3(G169gat), .A4(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n862_), .B1(new_n804_), .B2(new_n808_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n233_), .A2(new_n297_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT126), .Z(new_n869_));
  AND2_X1   g668(.A1(new_n863_), .A2(G169gat), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n864_), .B(KEYINPUT125), .Z(new_n871_));
  OAI221_X1 g670(.A(new_n866_), .B1(new_n867_), .B2(new_n869_), .C1(new_n870_), .C2(new_n871_), .ZN(G1348gat));
  INV_X1    g671(.A(new_n867_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G176gat), .B1(new_n873_), .B2(new_n602_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n435_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n861_), .A2(new_n246_), .A3(new_n523_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(G1349gat));
  NOR3_X1   g676(.A1(new_n867_), .A2(new_n265_), .A3(new_n538_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n875_), .A2(new_n288_), .A3(new_n539_), .A4(new_n860_), .ZN(new_n879_));
  INV_X1    g678(.A(G183gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(G1350gat));
  OAI21_X1  g680(.A(G190gat), .B1(new_n867_), .B2(new_n572_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n578_), .A2(new_n306_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n867_), .B2(new_n883_), .ZN(G1351gat));
  NAND4_X1  g683(.A1(new_n842_), .A2(new_n233_), .A3(new_n843_), .A4(new_n860_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g685(.A1(new_n842_), .A2(new_n602_), .A3(new_n843_), .A4(new_n860_), .ZN(new_n887_));
  INV_X1    g686(.A(G204gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n854_), .A2(new_n310_), .A3(new_n602_), .A4(new_n860_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1353gat));
  AOI21_X1  g690(.A(new_n538_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n842_), .A2(new_n843_), .A3(new_n860_), .A4(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT127), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n893_), .B(new_n895_), .ZN(G1354gat));
  INV_X1    g695(.A(G218gat), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n854_), .A2(new_n897_), .A3(new_n578_), .A4(new_n860_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n854_), .A2(new_n571_), .A3(new_n860_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1355gat));
endmodule


