//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n939_, new_n940_, new_n941_,
    new_n943_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_, new_n974_, new_n975_, new_n976_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n983_, new_n984_, new_n986_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n993_, new_n994_,
    new_n995_;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203_));
  XOR2_X1   g002(.A(G29gat), .B(G36gat), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT73), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G29gat), .B(G36gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT73), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n203_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n206_), .A2(new_n208_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n209_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(KEYINPUT15), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  INV_X1    g023(.A(G92gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT9), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT9), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(G85gat), .A3(G92gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n223_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n232_), .A2(KEYINPUT64), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT64), .B1(new_n232_), .B2(new_n233_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n231_), .B1(new_n236_), .B2(G106gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n238_));
  OR3_X1    g037(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n223_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT8), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n226_), .A2(new_n227_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n241_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n237_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n218_), .A2(KEYINPUT74), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT74), .B1(new_n218_), .B2(new_n245_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n202_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n215_), .A2(new_n216_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n251_));
  AND2_X1   g050(.A1(G232gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n253_), .A2(KEYINPUT35), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(KEYINPUT35), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT72), .Z(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n248_), .A2(new_n256_), .A3(new_n259_), .ZN(new_n260_));
  OAI221_X1 g059(.A(new_n255_), .B1(new_n202_), .B2(new_n258_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT77), .A3(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G190gat), .B(G218gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT76), .ZN(new_n264_));
  XOR2_X1   g063(.A(G134gat), .B(G162gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT36), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n262_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n268_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n260_), .A2(KEYINPUT77), .A3(new_n261_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT37), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n260_), .A2(new_n261_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n266_), .A2(new_n267_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n272_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT78), .B(G8gat), .ZN(new_n280_));
  INV_X1    g079(.A(G1gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT14), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G15gat), .B(G22gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G1gat), .B(G8gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G231gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT65), .B(G71gat), .ZN(new_n289_));
  INV_X1    g088(.A(G78gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(G71gat), .ZN(new_n293_));
  INV_X1    g092(.A(G71gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(KEYINPUT65), .ZN(new_n295_));
  OAI21_X1  g094(.A(G78gat), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G64gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G57gat), .ZN(new_n299_));
  INV_X1    g098(.A(G57gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G64gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n301_), .A3(KEYINPUT11), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n302_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT11), .B1(new_n299_), .B2(new_n301_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n296_), .B(new_n291_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n288_), .B(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G127gat), .B(G155gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G183gat), .B(G211gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT17), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n313_), .A2(KEYINPUT17), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n308_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n279_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT13), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT70), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G120gat), .B(G148gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT5), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G176gat), .B(G204gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT66), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n303_), .A2(new_n306_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n329_), .B1(new_n245_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n240_), .A2(new_n242_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT8), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n307_), .A2(new_n336_), .A3(KEYINPUT66), .A4(new_n237_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n331_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n332_), .B1(new_n331_), .B2(new_n337_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n307_), .B1(new_n237_), .B2(new_n336_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G230gat), .A2(G233gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n328_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n331_), .A2(new_n337_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT67), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n245_), .A2(new_n330_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n331_), .A2(new_n337_), .A3(new_n332_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n342_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT68), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n343_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n342_), .B1(new_n245_), .B2(new_n330_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n346_), .A2(KEYINPUT12), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT12), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n245_), .B2(new_n330_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n353_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT69), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n340_), .A2(new_n355_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n356_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(KEYINPUT69), .A3(new_n353_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n327_), .B1(new_n351_), .B2(new_n365_), .ZN(new_n366_));
  AOI211_X1 g165(.A(new_n326_), .B(new_n364_), .C1(new_n343_), .C2(new_n350_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n322_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n348_), .A2(KEYINPUT68), .A3(new_n349_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT68), .B1(new_n348_), .B2(new_n349_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n365_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n326_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n351_), .A2(new_n365_), .A3(new_n327_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n368_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n320_), .A2(new_n378_), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n379_), .A2(KEYINPUT80), .ZN(new_n380_));
  INV_X1    g179(.A(G169gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT22), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G169gat), .ZN(new_n384_));
  INV_X1    g183(.A(G176gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT22), .B(G169gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(KEYINPUT84), .A3(new_n385_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT23), .ZN(new_n394_));
  OR2_X1    g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n392_), .A2(KEYINPUT85), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT85), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n388_), .A2(new_n390_), .A3(new_n397_), .A4(new_n391_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT25), .B(G183gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G190gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT24), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G169gat), .A2(G176gat), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n399_), .A2(new_n400_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(KEYINPUT24), .A3(new_n391_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n394_), .A2(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n396_), .A2(new_n398_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408_));
  INV_X1    g207(.A(G15gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT30), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n392_), .A2(KEYINPUT85), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n394_), .A2(new_n395_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n398_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n403_), .A2(new_n394_), .A3(new_n405_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n411_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n412_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G134gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(G127gat), .ZN(new_n422_));
  INV_X1    g221(.A(G127gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(G134gat), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n422_), .A2(new_n424_), .A3(KEYINPUT86), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT86), .B1(new_n422_), .B2(new_n424_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G113gat), .B(G120gat), .Z(new_n427_));
  NOR3_X1   g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G113gat), .B(G120gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT86), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n423_), .A2(G134gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n421_), .A2(G127gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n422_), .A2(new_n424_), .A3(KEYINPUT86), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n429_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n428_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n420_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438_));
  INV_X1    g237(.A(G43gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT31), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n412_), .B(new_n419_), .C1(new_n428_), .C2(new_n435_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n437_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446_));
  INV_X1    g245(.A(G155gat), .ZN(new_n447_));
  INV_X1    g246(.A(G162gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT1), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G155gat), .A2(G162gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n446_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT1), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n453_), .B1(G155gat), .B2(G162gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(KEYINPUT88), .A3(new_n450_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n450_), .A2(KEYINPUT1), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n452_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  OR3_X1    g257(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n459_), .A2(new_n460_), .B1(G141gat), .B2(G148gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464_));
  INV_X1    g263(.A(G141gat), .ZN(new_n465_));
  INV_X1    g264(.A(G148gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT3), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT3), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n464_), .A2(new_n469_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT2), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n471_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n468_), .A2(new_n470_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G155gat), .A2(G162gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n451_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n462_), .A2(new_n463_), .A3(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(KEYINPUT28), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT28), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n458_), .A2(new_n461_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n481_), .B2(new_n463_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G22gat), .B(G50gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n479_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n478_), .A2(KEYINPUT28), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n481_), .A2(new_n480_), .A3(new_n463_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n483_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G228gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n463_), .B1(new_n462_), .B2(new_n477_), .ZN(new_n494_));
  OR2_X1    g293(.A1(G197gat), .A2(G204gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G197gat), .A2(G204gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(KEYINPUT21), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G211gat), .B(G218gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n499_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n495_), .A2(new_n496_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT21), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n497_), .A2(new_n498_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n501_), .A2(new_n502_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n493_), .B1(new_n494_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n505_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n502_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n509_), .B1(new_n510_), .B2(new_n500_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n511_), .B(new_n492_), .C1(new_n481_), .C2(new_n463_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n491_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n508_), .A2(new_n512_), .A3(new_n491_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n489_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT93), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n489_), .A2(new_n514_), .A3(new_n518_), .A4(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n515_), .B1(new_n513_), .B2(KEYINPUT91), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n508_), .A2(new_n523_), .A3(new_n512_), .A4(new_n491_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n489_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n521_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  AOI211_X1 g326(.A(KEYINPUT92), .B(new_n489_), .C1(new_n522_), .C2(new_n524_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n520_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n454_), .A2(KEYINPUT88), .A3(new_n450_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT88), .B1(new_n454_), .B2(new_n450_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n456_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n461_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n477_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT96), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n436_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT96), .B1(new_n428_), .B2(new_n435_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n427_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n433_), .A2(new_n434_), .A3(new_n429_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(new_n535_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n537_), .A2(new_n481_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G225gat), .A2(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT4), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT97), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n547_), .A2(new_n481_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT4), .B1(new_n538_), .B2(new_n539_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT97), .B1(new_n534_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n545_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n546_), .B1(new_n536_), .B2(new_n541_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT98), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT98), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n537_), .A2(new_n481_), .A3(new_n540_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n540_), .B1(new_n537_), .B2(new_n481_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT4), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n548_), .B1(new_n547_), .B2(new_n481_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n534_), .A2(KEYINPUT97), .A3(new_n550_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n543_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n555_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n544_), .B1(new_n554_), .B2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G1gat), .B(G29gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT100), .ZN(new_n565_));
  XOR2_X1   g364(.A(G57gat), .B(G85gat), .Z(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n567_), .A2(new_n570_), .A3(new_n568_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n563_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n544_), .A2(new_n574_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(new_n554_), .B2(new_n562_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT103), .B(KEYINPUT27), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n507_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G226gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT19), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n386_), .A2(new_n391_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n414_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n416_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT20), .B1(new_n511_), .B2(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n582_), .A2(new_n584_), .A3(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n584_), .B(KEYINPUT94), .Z(new_n590_));
  NAND3_X1  g389(.A1(new_n415_), .A2(new_n507_), .A3(new_n416_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT20), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n511_), .B2(new_n587_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n590_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G8gat), .B(G36gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G64gat), .B(G92gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n589_), .A2(new_n594_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n591_), .A2(new_n593_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n590_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n406_), .A2(new_n403_), .B1(new_n585_), .B2(new_n414_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n592_), .B1(new_n507_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n584_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n606_), .B(new_n607_), .C1(new_n407_), .C2(new_n507_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n601_), .B1(new_n604_), .B2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n581_), .B1(new_n600_), .B2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n604_), .A2(new_n608_), .A3(new_n601_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n602_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n606_), .B1(new_n407_), .B2(new_n507_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n612_), .A2(new_n590_), .B1(new_n613_), .B2(new_n584_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n611_), .B(KEYINPUT27), .C1(new_n614_), .C2(new_n601_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n576_), .A2(new_n579_), .A3(new_n610_), .A4(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n445_), .B1(new_n529_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n525_), .A2(new_n526_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT92), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n525_), .A2(new_n521_), .A3(new_n526_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n545_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n574_), .B1(new_n558_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n542_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n536_), .A2(new_n541_), .A3(KEYINPUT102), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n545_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n623_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n599_), .B1(new_n589_), .B2(new_n594_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n628_), .A2(new_n611_), .A3(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n579_), .A2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT98), .B1(new_n552_), .B2(new_n553_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n558_), .A2(new_n555_), .A3(new_n561_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n577_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n631_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n632_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n601_), .A2(KEYINPUT32), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n613_), .A2(new_n584_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n591_), .A2(new_n593_), .A3(new_n590_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n639_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n589_), .A2(new_n594_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n643_), .B2(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n633_), .A2(new_n634_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n574_), .B1(new_n645_), .B2(new_n544_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n644_), .B1(new_n646_), .B2(new_n635_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n621_), .A2(new_n638_), .A3(new_n647_), .A4(new_n520_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n617_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n617_), .B2(new_n648_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n646_), .A2(new_n635_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n445_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n610_), .A2(new_n615_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n653_), .A2(new_n529_), .A3(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n650_), .A2(new_n651_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n218_), .A2(new_n286_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT81), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n218_), .A2(KEYINPUT81), .A3(new_n286_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n286_), .A2(new_n249_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(G229gat), .A2(G233gat), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n286_), .B(new_n249_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT83), .ZN(new_n670_));
  XOR2_X1   g469(.A(G113gat), .B(G141gat), .Z(new_n671_));
  XNOR2_X1  g470(.A(G169gat), .B(G197gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT82), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n669_), .A2(new_n670_), .A3(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n665_), .A2(new_n668_), .A3(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n670_), .B1(new_n669_), .B2(new_n675_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n656_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n379_), .A2(KEYINPUT80), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n380_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n652_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n380_), .A2(KEYINPUT105), .A3(new_n681_), .A4(new_n682_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n685_), .A2(new_n281_), .A3(new_n686_), .A4(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT38), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n689_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n680_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT106), .B1(new_n377_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  AOI211_X1 g493(.A(new_n694_), .B(new_n680_), .C1(new_n368_), .C2(new_n376_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n272_), .A2(new_n276_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n617_), .A2(new_n648_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n655_), .B1(new_n698_), .B2(KEYINPUT104), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n617_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n696_), .A2(new_n319_), .A3(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT107), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(new_n686_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n690_), .B(new_n691_), .C1(new_n281_), .C2(new_n704_), .ZN(G1324gat));
  NAND4_X1  g504(.A1(new_n685_), .A2(new_n654_), .A3(new_n280_), .A4(new_n687_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n696_), .A2(new_n654_), .A3(new_n319_), .A4(new_n701_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G8gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT108), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT39), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n707_), .A2(new_n711_), .A3(G8gat), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n709_), .A2(new_n710_), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n709_), .B2(new_n712_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n706_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT40), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n706_), .B(KEYINPUT40), .C1(new_n713_), .C2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1325gat));
  INV_X1    g518(.A(new_n683_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n409_), .A3(new_n445_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n409_), .B1(new_n703_), .B2(new_n445_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(KEYINPUT41), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(KEYINPUT41), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(G1326gat));
  INV_X1    g524(.A(G22gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(new_n726_), .A3(new_n529_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n703_), .B2(new_n529_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n729_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1327gat));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n697_), .A2(new_n733_), .A3(new_n318_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n269_), .A2(new_n271_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT110), .B1(new_n735_), .B2(new_n319_), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n734_), .A2(new_n736_), .B1(new_n368_), .B2(new_n376_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n681_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G29gat), .B1(new_n738_), .B2(new_n686_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n693_), .A2(new_n695_), .A3(new_n319_), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT43), .B(new_n279_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n698_), .A2(KEYINPUT104), .ZN(new_n743_));
  INV_X1    g542(.A(new_n655_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n700_), .A3(new_n744_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n277_), .A2(new_n278_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(KEYINPUT44), .B(new_n740_), .C1(new_n741_), .C2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n366_), .A2(new_n367_), .A3(new_n374_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n372_), .A2(new_n373_), .B1(KEYINPUT70), .B2(new_n321_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n692_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n694_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n377_), .A2(KEYINPUT106), .A3(new_n692_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n318_), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n656_), .B2(new_n279_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n745_), .A2(new_n742_), .A3(new_n746_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT109), .B1(new_n758_), .B2(KEYINPUT44), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n740_), .B1(new_n741_), .B2(new_n747_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n749_), .B1(new_n759_), .B2(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n686_), .A2(G29gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n739_), .B1(new_n764_), .B2(new_n765_), .ZN(G1328gat));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n748_), .A2(new_n654_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n758_), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n761_), .B1(new_n760_), .B2(new_n762_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(KEYINPUT112), .A2(G36gat), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G36gat), .B1(new_n610_), .B2(new_n615_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n745_), .A2(new_n737_), .A3(new_n692_), .A4(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT111), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n776_), .A2(KEYINPUT111), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n776_), .A2(KEYINPUT111), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(KEYINPUT45), .A3(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(KEYINPUT112), .A3(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n767_), .B1(new_n774_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n748_), .A2(new_n654_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n759_), .B2(new_n763_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n767_), .B(new_n783_), .C1(new_n786_), .C2(new_n772_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n784_), .A2(new_n788_), .ZN(G1329gat));
  AOI21_X1  g588(.A(G43gat), .B1(new_n738_), .B2(new_n445_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n445_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(new_n439_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n764_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT47), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n792_), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n796_), .B(new_n749_), .C1(new_n759_), .C2(new_n763_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT47), .B1(new_n797_), .B2(new_n790_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n795_), .A2(new_n798_), .ZN(G1330gat));
  AOI21_X1  g598(.A(G50gat), .B1(new_n738_), .B2(new_n529_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n529_), .ZN(new_n801_));
  INV_X1    g600(.A(G50gat), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n800_), .B1(new_n764_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n803_), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n807_), .B(new_n749_), .C1(new_n759_), .C2(new_n763_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT113), .B1(new_n808_), .B2(new_n800_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n809_), .ZN(G1331gat));
  NOR3_X1   g609(.A1(new_n377_), .A2(new_n692_), .A3(new_n318_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n701_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n701_), .A2(KEYINPUT114), .A3(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G57gat), .B1(new_n816_), .B2(new_n652_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n656_), .A2(new_n692_), .A3(new_n377_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n320_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n300_), .A3(new_n686_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n821_), .ZN(G1332gat));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n298_), .A3(new_n654_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n816_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n654_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n826_));
  AND3_X1   g625(.A1(new_n825_), .A2(G64gat), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n825_), .B2(G64gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n823_), .B1(new_n827_), .B2(new_n828_), .ZN(G1333gat));
  NAND3_X1  g628(.A1(new_n820_), .A2(new_n294_), .A3(new_n445_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n814_), .A2(new_n445_), .A3(new_n815_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n831_), .A2(new_n832_), .A3(G71gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n831_), .B2(G71gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n830_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1334gat));
  NAND3_X1  g636(.A1(new_n820_), .A2(new_n290_), .A3(new_n529_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G78gat), .B1(new_n816_), .B2(new_n801_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n839_), .A2(KEYINPUT50), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(KEYINPUT50), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n838_), .B1(new_n840_), .B2(new_n841_), .ZN(G1335gat));
  AND2_X1   g641(.A1(new_n734_), .A2(new_n736_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n818_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n224_), .B1(new_n845_), .B2(new_n652_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n756_), .A2(new_n757_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n377_), .A2(new_n692_), .A3(new_n319_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n686_), .A2(G85gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT117), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n846_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT118), .ZN(G1336gat));
  AOI21_X1  g652(.A(new_n849_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n654_), .A2(new_n225_), .ZN(new_n855_));
  OAI22_X1  g654(.A1(new_n854_), .A2(new_n225_), .B1(new_n845_), .B2(new_n855_), .ZN(G1337gat));
  NOR2_X1   g655(.A1(new_n791_), .A2(new_n236_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n818_), .A2(new_n844_), .A3(new_n857_), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(KEYINPUT119), .Z(new_n859_));
  OAI21_X1  g658(.A(G99gat), .B1(new_n849_), .B2(new_n791_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g661(.A1(new_n845_), .A2(G106gat), .A3(new_n801_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n847_), .A2(new_n529_), .A3(new_n848_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n864_), .A2(new_n865_), .A3(G106gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n864_), .B2(G106gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n863_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n362_), .A2(new_n331_), .A3(new_n337_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n352_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n871_), .A2(new_n349_), .B1(new_n872_), .B2(KEYINPUT55), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n359_), .A2(new_n363_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n327_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n876_), .A2(KEYINPUT56), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(KEYINPUT56), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n680_), .A2(new_n367_), .ZN(new_n881_));
  OR3_X1    g680(.A1(new_n876_), .A2(new_n878_), .A3(KEYINPUT56), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n661_), .A2(new_n662_), .A3(new_n667_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n673_), .B1(new_n666_), .B2(new_n663_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n677_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n883_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n870_), .B1(new_n889_), .B2(new_n697_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n697_), .B1(new_n883_), .B2(new_n888_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT57), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n877_), .A2(new_n879_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n373_), .A2(new_n887_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n893_), .B(new_n894_), .C1(KEYINPUT122), .C2(KEYINPUT58), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(new_n746_), .A3(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n890_), .A2(new_n892_), .A3(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n819_), .A2(new_n680_), .A3(new_n377_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n379_), .B(new_n680_), .C1(KEYINPUT120), .C2(new_n904_), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n900_), .A2(new_n318_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n529_), .A2(new_n654_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(new_n686_), .A3(new_n445_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT59), .B1(new_n906_), .B2(new_n908_), .ZN(new_n909_));
  AOI211_X1 g708(.A(new_n870_), .B(new_n697_), .C1(new_n883_), .C2(new_n888_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n899_), .B1(new_n891_), .B2(KEYINPUT57), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(KEYINPUT123), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n890_), .A2(new_n913_), .A3(new_n899_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n319_), .B1(new_n912_), .B2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n903_), .A2(new_n905_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n908_), .A2(KEYINPUT59), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n909_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(G113gat), .B1(new_n920_), .B2(new_n680_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n906_), .A2(new_n908_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  OR3_X1    g722(.A1(new_n923_), .A2(G113gat), .A3(new_n680_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n921_), .A2(new_n924_), .ZN(G1340gat));
  OAI21_X1  g724(.A(G120gat), .B1(new_n920_), .B2(new_n377_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n377_), .A2(KEYINPUT60), .ZN(new_n927_));
  MUX2_X1   g726(.A(new_n927_), .B(KEYINPUT60), .S(G120gat), .Z(new_n928_));
  NAND2_X1  g727(.A1(new_n922_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n929_), .ZN(G1341gat));
  OAI21_X1  g729(.A(new_n423_), .B1(new_n923_), .B2(new_n318_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n318_), .A2(new_n423_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT124), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n909_), .B(new_n933_), .C1(new_n918_), .C2(new_n919_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n931_), .A2(new_n934_), .ZN(G1342gat));
  OAI21_X1  g734(.A(G134gat), .B1(new_n920_), .B2(new_n279_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n922_), .A2(new_n421_), .A3(new_n697_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1343gat));
  NOR2_X1   g737(.A1(new_n906_), .A2(new_n445_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n801_), .A2(new_n652_), .A3(new_n654_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n939_), .A2(new_n692_), .A3(new_n940_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g741(.A1(new_n939_), .A2(new_n378_), .A3(new_n940_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g743(.A1(new_n939_), .A2(new_n319_), .A3(new_n940_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(KEYINPUT61), .B(G155gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(G1346gat));
  AND4_X1   g746(.A1(G162gat), .A2(new_n939_), .A3(new_n746_), .A4(new_n940_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n318_), .B1(new_n911_), .B2(new_n910_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n916_), .A2(new_n949_), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n950_), .A2(new_n791_), .A3(new_n697_), .A4(new_n940_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(new_n448_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(KEYINPUT125), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n951_), .A2(new_n954_), .A3(new_n448_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n948_), .B1(new_n953_), .B2(new_n955_), .ZN(G1347gat));
  NAND2_X1  g755(.A1(new_n652_), .A2(new_n654_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n957_), .A2(new_n791_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n959_), .A2(new_n529_), .ZN(new_n960_));
  OAI211_X1 g759(.A(new_n692_), .B(new_n960_), .C1(new_n915_), .C2(new_n917_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(G169gat), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  INV_X1    g763(.A(new_n960_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n918_), .A2(new_n965_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n966_), .A2(new_n389_), .A3(new_n692_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n961_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n964_), .A2(new_n967_), .A3(new_n968_), .ZN(G1348gat));
  NAND2_X1  g768(.A1(new_n966_), .A2(new_n378_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n906_), .A2(new_n529_), .ZN(new_n971_));
  NOR3_X1   g770(.A1(new_n377_), .A2(new_n385_), .A3(new_n959_), .ZN(new_n972_));
  AOI22_X1  g771(.A1(new_n970_), .A2(new_n385_), .B1(new_n971_), .B2(new_n972_), .ZN(G1349gat));
  NOR2_X1   g772(.A1(new_n959_), .A2(new_n318_), .ZN(new_n974_));
  AOI21_X1  g773(.A(G183gat), .B1(new_n971_), .B2(new_n974_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n318_), .A2(new_n399_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n975_), .B1(new_n966_), .B2(new_n976_), .ZN(G1350gat));
  NAND3_X1  g776(.A1(new_n966_), .A2(new_n400_), .A3(new_n697_), .ZN(new_n978_));
  OAI211_X1 g777(.A(new_n746_), .B(new_n960_), .C1(new_n915_), .C2(new_n917_), .ZN(new_n979_));
  AND3_X1   g778(.A1(new_n979_), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n980_));
  AOI21_X1  g779(.A(KEYINPUT126), .B1(new_n979_), .B2(G190gat), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n978_), .B1(new_n980_), .B2(new_n981_), .ZN(G1351gat));
  NOR2_X1   g781(.A1(new_n801_), .A2(new_n957_), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n939_), .A2(new_n692_), .A3(new_n983_), .ZN(new_n984_));
  XNOR2_X1  g783(.A(new_n984_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g784(.A1(new_n939_), .A2(new_n378_), .A3(new_n983_), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n986_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g786(.A(new_n318_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(KEYINPUT127), .ZN(new_n989_));
  NAND3_X1  g788(.A1(new_n939_), .A2(new_n983_), .A3(new_n989_), .ZN(new_n990_));
  OR2_X1    g789(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n991_));
  XNOR2_X1  g790(.A(new_n990_), .B(new_n991_), .ZN(G1354gat));
  NAND2_X1  g791(.A1(new_n939_), .A2(new_n983_), .ZN(new_n993_));
  OAI21_X1  g792(.A(G218gat), .B1(new_n993_), .B2(new_n279_), .ZN(new_n994_));
  OR2_X1    g793(.A1(new_n735_), .A2(G218gat), .ZN(new_n995_));
  OAI21_X1  g794(.A(new_n994_), .B1(new_n993_), .B2(new_n995_), .ZN(G1355gat));
endmodule


