//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n583_, new_n584_, new_n585_, new_n586_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n819_, new_n820_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(new_n202_), .A2(KEYINPUT74), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(KEYINPUT74), .ZN(new_n204_));
  XOR2_X1   g003(.A(G43gat), .B(G50gat), .Z(new_n205_));
  OR3_X1    g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT78), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210_));
  INV_X1    g009(.A(G1gat), .ZN(new_n211_));
  INV_X1    g010(.A(G8gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G1gat), .B(G8gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n214_), .B(new_n215_), .Z(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n209_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n209_), .A2(new_n217_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G229gat), .A3(G233gat), .ZN(new_n221_));
  XOR2_X1   g020(.A(new_n208_), .B(KEYINPUT15), .Z(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n217_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n218_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G141gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G169gat), .B(G197gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT79), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n231_), .B(KEYINPUT80), .Z(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n226_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n221_), .A2(new_n232_), .A3(new_n225_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT104), .B(KEYINPUT27), .Z(new_n237_));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT84), .B1(new_n238_), .B2(KEYINPUT23), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(KEYINPUT23), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  NOR3_X1   g040(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n242_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT25), .B(G183gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT26), .B(G190gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n241_), .A2(new_n246_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(KEYINPUT82), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n238_), .A2(KEYINPUT23), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n238_), .B2(KEYINPUT23), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(G183gat), .B2(G190gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT98), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n245_), .B(KEYINPUT96), .Z(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT22), .B(G169gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT97), .Z(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n260_), .B2(G176gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n250_), .B1(new_n257_), .B2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT91), .B(G197gat), .Z(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(G204gat), .ZN(new_n265_));
  INV_X1    g064(.A(G197gat), .ZN(new_n266_));
  INV_X1    g065(.A(G204gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT21), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G197gat), .A2(G204gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n264_), .B2(G204gat), .ZN(new_n271_));
  OAI221_X1 g070(.A(new_n263_), .B1(new_n265_), .B2(new_n268_), .C1(new_n269_), .C2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G211gat), .B(G218gat), .Z(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(KEYINPUT21), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n262_), .A2(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(KEYINPUT93), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT81), .B(G190gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n241_), .B1(G183gat), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT83), .B(G169gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n278_), .B2(KEYINPUT26), .ZN(new_n285_));
  INV_X1    g084(.A(new_n247_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n255_), .B(new_n246_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n275_), .A2(KEYINPUT93), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n277_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT19), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT20), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n276_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n288_), .B1(new_n277_), .B2(new_n289_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n262_), .A2(new_n275_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(KEYINPUT99), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(KEYINPUT99), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n295_), .B1(new_n301_), .B2(new_n292_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G8gat), .B(G36gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT18), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G64gat), .B(G92gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  NOR2_X1   g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n306_), .ZN(new_n308_));
  AOI211_X1 g107(.A(new_n308_), .B(new_n295_), .C1(new_n301_), .C2(new_n292_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n237_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n311_));
  NAND3_X1  g110(.A1(new_n276_), .A2(new_n290_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n292_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(new_n301_), .B2(new_n292_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n306_), .B(KEYINPUT103), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n302_), .A2(new_n306_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(KEYINPUT27), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n310_), .A2(new_n318_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT3), .ZN(new_n321_));
  INV_X1    g120(.A(G141gat), .ZN(new_n322_));
  INV_X1    g121(.A(G148gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324_));
  OAI22_X1  g123(.A1(new_n322_), .A2(new_n323_), .B1(new_n324_), .B2(KEYINPUT87), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(KEYINPUT2), .ZN(new_n327_));
  OAI211_X1 g126(.A(KEYINPUT87), .B(new_n324_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n321_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT88), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n330_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n333_), .B(KEYINPUT89), .Z(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G141gat), .B(G148gat), .Z(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n336_), .B(new_n337_), .C1(KEYINPUT1), .C2(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n340_));
  OR3_X1    g139(.A1(new_n339_), .A2(KEYINPUT29), .A3(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G22gat), .B(G50gat), .Z(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n339_), .B2(KEYINPUT29), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n342_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n339_), .A2(KEYINPUT29), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n275_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(G228gat), .A3(G233gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G228gat), .A2(G233gat), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n347_), .A2(new_n350_), .A3(new_n289_), .A4(new_n277_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n353_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n346_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT94), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT94), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n346_), .B(new_n359_), .C1(new_n354_), .C2(new_n356_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n346_), .A2(new_n356_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n349_), .A2(new_n351_), .A3(KEYINPUT95), .A4(new_n355_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT95), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n358_), .A2(new_n360_), .A3(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n319_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(G43gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n288_), .B(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  INV_X1    g172(.A(G15gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT30), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G127gat), .B(G134gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  XNOR2_X1  g178(.A(new_n376_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n372_), .B(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n335_), .A2(new_n338_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n379_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT100), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n339_), .B2(new_n379_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n382_), .A2(new_n385_), .A3(new_n383_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT4), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n384_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(G85gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT0), .B(G57gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n384_), .A2(new_n386_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n388_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n393_), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n395_), .A2(new_n400_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n393_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n403_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n399_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT102), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n395_), .A2(KEYINPUT102), .A3(new_n400_), .A4(new_n403_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n381_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n367_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT105), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT105), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n367_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n314_), .A2(KEYINPUT32), .A3(new_n306_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n306_), .A2(KEYINPUT32), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n302_), .A2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n409_), .A2(new_n410_), .A3(new_n417_), .A4(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n407_), .A2(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(KEYINPUT33), .B(new_n399_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n307_), .A2(new_n309_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n401_), .A2(new_n402_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n399_), .B1(new_n425_), .B2(new_n394_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .A4(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n366_), .B1(new_n420_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n409_), .A2(new_n410_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n310_), .A2(new_n318_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n366_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n381_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n236_), .B1(new_n416_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT8), .ZN(new_n436_));
  XOR2_X1   g235(.A(G85gat), .B(G92gat), .Z(new_n437_));
  NAND2_X1  g236(.A1(G99gat), .A2(G106gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT7), .ZN(new_n441_));
  INV_X1    g240(.A(G99gat), .ZN(new_n442_));
  INV_X1    g241(.A(G106gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n436_), .B(new_n437_), .C1(new_n440_), .C2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT69), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(KEYINPUT6), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n439_), .A2(KEYINPUT67), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n438_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT68), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n444_), .A2(new_n453_), .A3(new_n445_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n439_), .A2(KEYINPUT67), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(KEYINPUT6), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(G99gat), .A4(G106gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n452_), .A2(new_n454_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n453_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n448_), .B(new_n437_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT8), .ZN(new_n461_));
  INV_X1    g260(.A(new_n459_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(new_n454_), .A3(new_n452_), .A4(new_n457_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n448_), .B1(new_n463_), .B2(new_n437_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n447_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT66), .B(G92gat), .ZN(new_n466_));
  INV_X1    g265(.A(G85gat), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n466_), .A2(KEYINPUT9), .A3(new_n467_), .ZN(new_n468_));
  AOI211_X1 g267(.A(new_n440_), .B(new_n468_), .C1(KEYINPUT9), .C2(new_n437_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT10), .B(G99gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT64), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n472_), .A2(KEYINPUT65), .A3(new_n443_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT65), .B1(new_n472_), .B2(new_n443_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n469_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n465_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G57gat), .B(G64gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n478_));
  XOR2_X1   g277(.A(G71gat), .B(G78gat), .Z(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n479_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n476_), .A2(KEYINPUT12), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT70), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n465_), .A2(new_n487_), .A3(new_n475_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n487_), .B1(new_n465_), .B2(new_n475_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n484_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT12), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n486_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(G230gat), .ZN(new_n493_));
  INV_X1    g292(.A(G233gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n488_), .A2(new_n489_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(new_n483_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n476_), .A2(KEYINPUT70), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n465_), .A2(new_n487_), .A3(new_n475_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n483_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n490_), .A2(new_n500_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n492_), .A2(new_n497_), .B1(new_n501_), .B2(new_n495_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G120gat), .B(G148gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G176gat), .B(G204gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n502_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT72), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n502_), .A2(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n510_), .A2(new_n511_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n515_));
  OAI22_X1  g314(.A1(new_n513_), .A2(new_n514_), .B1(KEYINPUT73), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n514_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n512_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT35), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT34), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n496_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n222_), .A2(new_n476_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n527_));
  AOI211_X1 g326(.A(new_n522_), .B(new_n525_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n527_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n525_), .A2(new_n522_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G190gat), .B(G218gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT75), .ZN(new_n534_));
  XOR2_X1   g333(.A(G134gat), .B(G162gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n532_), .A2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n536_), .A2(new_n537_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n538_), .B(new_n541_), .C1(new_n531_), .C2(new_n528_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n544_));
  NAND2_X1  g343(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n540_), .A2(KEYINPUT76), .A3(new_n542_), .A4(KEYINPUT37), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n216_), .B(new_n483_), .Z(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G127gat), .B(G155gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT16), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G183gat), .B(G211gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n551_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n555_), .A2(new_n556_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n558_), .B1(new_n559_), .B2(new_n551_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT77), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n548_), .A2(new_n561_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n435_), .A2(new_n521_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n430_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n211_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT38), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n563_), .A2(KEYINPUT38), .A3(new_n211_), .A4(new_n564_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n543_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n416_), .B2(new_n433_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n561_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n521_), .A2(new_n236_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(G1gat), .B1(new_n573_), .B2(new_n430_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n567_), .A2(new_n568_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT106), .ZN(G1324gat));
  NAND3_X1  g375(.A1(new_n563_), .A2(new_n212_), .A3(new_n319_), .ZN(new_n577_));
  OAI21_X1  g376(.A(G8gat), .B1(new_n573_), .B2(new_n431_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n578_), .A2(KEYINPUT39), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(KEYINPUT39), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n577_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g381(.A(G15gat), .B1(new_n573_), .B2(new_n381_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT41), .Z(new_n584_));
  INV_X1    g383(.A(new_n381_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n563_), .A2(new_n374_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(G1326gat));
  INV_X1    g386(.A(G22gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n573_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n589_), .B2(new_n366_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT42), .Z(new_n591_));
  NAND2_X1  g390(.A1(new_n366_), .A2(new_n588_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT107), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n563_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(G1327gat));
  INV_X1    g394(.A(new_n236_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n520_), .A2(new_n596_), .A3(new_n571_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT43), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n416_), .A2(new_n433_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n548_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT43), .B(new_n548_), .C1(new_n416_), .C2(new_n433_), .ZN(new_n603_));
  OAI211_X1 g402(.A(KEYINPUT44), .B(new_n598_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT43), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n600_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n597_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n604_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G29gat), .B1(new_n610_), .B2(new_n430_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n543_), .A2(new_n561_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n521_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n434_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n430_), .A2(G29gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT109), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n611_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT110), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT110), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(new_n622_), .A3(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(G1328gat));
  INV_X1    g423(.A(KEYINPUT46), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT112), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n431_), .A2(G36gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n434_), .A2(new_n614_), .A3(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n628_), .A2(KEYINPUT45), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(KEYINPUT45), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n604_), .B(new_n319_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(G36gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT112), .B1(new_n625_), .B2(KEYINPUT111), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1329gat));
  NAND2_X1  g434(.A1(new_n585_), .A2(G43gat), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n615_), .A2(new_n381_), .ZN(new_n637_));
  OAI22_X1  g436(.A1(new_n610_), .A2(new_n636_), .B1(G43gat), .B2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g438(.A(G50gat), .B1(new_n616_), .B2(new_n366_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n610_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n366_), .A2(G50gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n640_), .B1(new_n641_), .B2(new_n642_), .ZN(G1331gat));
  INV_X1    g442(.A(KEYINPUT113), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n600_), .B2(new_n236_), .ZN(new_n645_));
  AOI211_X1 g444(.A(KEYINPUT113), .B(new_n596_), .C1(new_n416_), .C2(new_n433_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n647_), .A2(new_n520_), .A3(new_n562_), .ZN(new_n648_));
  INV_X1    g447(.A(G57gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n564_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n520_), .A2(new_n596_), .A3(new_n571_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n570_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G57gat), .B1(new_n652_), .B2(new_n430_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(G1332gat));
  INV_X1    g453(.A(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n319_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G64gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT114), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT114), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n659_), .A3(G64gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n658_), .A2(KEYINPUT48), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(G64gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n648_), .A2(new_n662_), .A3(new_n319_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT48), .B1(new_n658_), .B2(new_n660_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1333gat));
  NOR2_X1   g465(.A1(new_n381_), .A2(G71gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT115), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n648_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G71gat), .B1(new_n652_), .B2(new_n381_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(KEYINPUT49), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(KEYINPUT49), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n669_), .B1(new_n671_), .B2(new_n672_), .ZN(G1334gat));
  INV_X1    g472(.A(G78gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n648_), .A2(new_n674_), .A3(new_n366_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n655_), .A2(new_n366_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G78gat), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT50), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT50), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(G1335gat));
  INV_X1    g479(.A(new_n647_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n520_), .A2(new_n613_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n681_), .A2(new_n467_), .A3(new_n564_), .A4(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT117), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT116), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n606_), .A2(new_n607_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n520_), .A2(new_n596_), .A3(new_n561_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(KEYINPUT116), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n684_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n686_), .A2(new_n685_), .A3(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(KEYINPUT116), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(KEYINPUT117), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n691_), .A2(new_n564_), .A3(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n683_), .B1(new_n695_), .B2(new_n467_), .ZN(G1336gat));
  AND2_X1   g495(.A1(new_n691_), .A2(new_n694_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n431_), .A2(new_n466_), .ZN(new_n698_));
  INV_X1    g497(.A(G92gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n681_), .A2(new_n319_), .A3(new_n682_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n697_), .A2(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(G1337gat));
  AND2_X1   g500(.A1(new_n585_), .A2(new_n472_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n682_), .B(new_n702_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT118), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n381_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n442_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT51), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT51), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n705_), .B(new_n709_), .C1(new_n706_), .C2(new_n442_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1338gat));
  NAND4_X1  g510(.A1(new_n681_), .A2(new_n443_), .A3(new_n366_), .A4(new_n682_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n366_), .B(new_n687_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT52), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G106gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G106gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g517(.A1(new_n561_), .A2(KEYINPUT119), .A3(new_n236_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT119), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(new_n571_), .B2(new_n596_), .ZN(new_n721_));
  AND4_X1   g520(.A1(new_n546_), .A2(new_n547_), .A3(new_n719_), .A4(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT54), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n520_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n722_), .B2(new_n520_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n596_), .A2(new_n509_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT120), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n483_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n500_), .B(new_n485_), .C1(new_n729_), .C2(KEYINPUT12), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n485_), .B1(new_n729_), .B2(KEYINPUT12), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n500_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT55), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n492_), .A2(new_n734_), .A3(new_n497_), .ZN(new_n735_));
  AOI221_X4 g534(.A(new_n728_), .B1(new_n495_), .B2(new_n730_), .C1(new_n733_), .C2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n735_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n730_), .A2(new_n495_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT120), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n507_), .B1(new_n736_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT56), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n492_), .A2(new_n734_), .A3(new_n497_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n734_), .B1(new_n492_), .B2(new_n497_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n738_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n728_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n737_), .A2(KEYINPUT120), .A3(new_n738_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(KEYINPUT56), .A3(new_n507_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n727_), .B1(new_n742_), .B2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n226_), .A2(new_n229_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n218_), .A2(new_n219_), .A3(new_n224_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n218_), .A2(new_n223_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT121), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n754_), .B2(new_n224_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n751_), .B1(new_n755_), .B2(new_n229_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n517_), .A2(new_n512_), .A3(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n543_), .B1(new_n750_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI211_X1 g559(.A(KEYINPUT57), .B(new_n543_), .C1(new_n750_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n756_), .A2(new_n509_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT56), .B1(new_n748_), .B2(new_n507_), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n741_), .B(new_n508_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT58), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT58), .B(new_n763_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n601_), .A3(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n760_), .A2(new_n761_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n726_), .B1(new_n771_), .B2(new_n571_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n564_), .A2(new_n367_), .A3(new_n585_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(G113gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n596_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n773_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n762_), .B1(new_n742_), .B2(new_n749_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n548_), .B1(new_n778_), .B2(KEYINPUT58), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n759_), .A2(new_n758_), .B1(new_n779_), .B2(new_n768_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n561_), .B1(new_n780_), .B2(new_n761_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT59), .B(new_n777_), .C1(new_n781_), .C2(new_n726_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT59), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n236_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n776_), .B1(new_n785_), .B2(new_n775_), .ZN(G1340gat));
  INV_X1    g585(.A(G120gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n520_), .B2(KEYINPUT60), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n774_), .B(new_n788_), .C1(KEYINPUT60), .C2(new_n787_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n520_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT122), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G120gat), .B1(new_n790_), .B2(new_n791_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(G1341gat));
  INV_X1    g593(.A(G127gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n774_), .A2(new_n795_), .A3(new_n561_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n571_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n795_), .ZN(G1342gat));
  INV_X1    g597(.A(G134gat), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n782_), .A2(new_n784_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n601_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n774_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n569_), .A2(new_n799_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT123), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT123), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n548_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n807_));
  OAI221_X1 g606(.A(new_n806_), .B1(new_n802_), .B2(new_n803_), .C1(new_n807_), .C2(new_n799_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n808_), .ZN(G1343gat));
  INV_X1    g608(.A(new_n772_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n366_), .A2(new_n381_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n811_), .A2(new_n430_), .A3(new_n319_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n236_), .ZN(new_n814_));
  XOR2_X1   g613(.A(KEYINPUT124), .B(G141gat), .Z(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(G1344gat));
  NOR2_X1   g615(.A1(new_n813_), .A2(new_n520_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(new_n323_), .ZN(G1345gat));
  NOR2_X1   g617(.A1(new_n813_), .A2(new_n571_), .ZN(new_n819_));
  XOR2_X1   g618(.A(KEYINPUT61), .B(G155gat), .Z(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1346gat));
  OAI21_X1  g620(.A(G162gat), .B1(new_n813_), .B2(new_n548_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n543_), .A2(G162gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n813_), .B2(new_n823_), .ZN(G1347gat));
  INV_X1    g623(.A(new_n411_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n825_), .A2(new_n366_), .A3(new_n431_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n772_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n596_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT62), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n829_), .A2(new_n830_), .A3(G169gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n829_), .B2(G169gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT125), .B1(new_n772_), .B2(new_n827_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n772_), .A2(KEYINPUT125), .A3(new_n827_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n236_), .A2(new_n260_), .ZN(new_n837_));
  OAI22_X1  g636(.A1(new_n831_), .A2(new_n832_), .B1(new_n836_), .B2(new_n837_), .ZN(G1348gat));
  INV_X1    g637(.A(new_n828_), .ZN(new_n839_));
  OAI21_X1  g638(.A(G176gat), .B1(new_n839_), .B2(new_n520_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n520_), .A2(G176gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n836_), .B2(new_n841_), .ZN(G1349gat));
  NAND2_X1  g641(.A1(new_n561_), .A2(new_n286_), .ZN(new_n843_));
  OR3_X1    g642(.A1(new_n772_), .A2(KEYINPUT125), .A3(new_n827_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n833_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n839_), .A2(new_n571_), .ZN(new_n846_));
  OAI22_X1  g645(.A1(new_n845_), .A2(KEYINPUT126), .B1(new_n846_), .B2(G183gat), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT126), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n836_), .A2(new_n848_), .A3(new_n843_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1350gat));
  OAI21_X1  g649(.A(G190gat), .B1(new_n836_), .B2(new_n548_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n569_), .A2(new_n248_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n836_), .B2(new_n852_), .ZN(G1351gat));
  NOR3_X1   g652(.A1(new_n564_), .A2(new_n431_), .A3(new_n811_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n810_), .A2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n236_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(new_n266_), .ZN(G1352gat));
  NOR2_X1   g656(.A1(new_n855_), .A2(new_n520_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n267_), .ZN(G1353gat));
  INV_X1    g658(.A(new_n855_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n571_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT127), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n862_), .B(new_n865_), .ZN(G1354gat));
  OR3_X1    g665(.A1(new_n855_), .A2(G218gat), .A3(new_n543_), .ZN(new_n867_));
  OAI21_X1  g666(.A(G218gat), .B1(new_n855_), .B2(new_n548_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1355gat));
endmodule


