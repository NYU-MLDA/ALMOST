//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT69), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n203_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT74), .B(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(KEYINPUT75), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(KEYINPUT75), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n206_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n213_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n214_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n203_), .B(new_n204_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(new_n215_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(new_n215_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(new_n206_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(KEYINPUT15), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT15), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n206_), .A2(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n221_), .A2(new_n229_), .A3(new_n231_), .A4(new_n215_), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n224_), .A2(new_n226_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G141gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G169gat), .B(G197gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT78), .B1(new_n233_), .B2(new_n236_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n216_), .A2(new_n206_), .A3(new_n217_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n222_), .B1(new_n221_), .B2(new_n215_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n226_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n232_), .A2(new_n218_), .A3(new_n225_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT78), .ZN(new_n243_));
  INV_X1    g042(.A(new_n236_), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT77), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n247_));
  AOI211_X1 g046(.A(KEYINPUT77), .B(new_n236_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n248_));
  OAI22_X1  g047(.A1(new_n237_), .A2(new_n245_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT96), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT19), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT87), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT22), .B(G169gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT89), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT79), .B(G176gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT90), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G183gat), .A2(G190gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT23), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(G183gat), .B2(G190gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT25), .B(G183gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(G190gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(KEYINPUT24), .A3(new_n260_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT88), .ZN(new_n275_));
  INV_X1    g074(.A(new_n265_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT24), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n276_), .B1(new_n277_), .B2(new_n271_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(KEYINPUT88), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n267_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT85), .B(G197gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G204gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(G197gat), .B2(G204gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G211gat), .B(G218gat), .Z(new_n287_));
  OR2_X1    g086(.A1(new_n282_), .A2(G204gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n285_), .B1(G197gat), .B2(G204gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT86), .ZN(new_n292_));
  INV_X1    g091(.A(new_n284_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(KEYINPUT21), .A3(new_n287_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n281_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT91), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT20), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n278_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n258_), .A2(new_n255_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n266_), .A2(new_n260_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n299_), .B1(new_n295_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n254_), .B1(new_n298_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G8gat), .B(G36gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT18), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G64gat), .B(G92gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  INV_X1    g110(.A(new_n295_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n299_), .B1(new_n312_), .B2(new_n303_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n253_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n281_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n313_), .B(new_n314_), .C1(new_n315_), .C2(new_n312_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n307_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT27), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n298_), .A2(new_n306_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n254_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n312_), .B1(new_n315_), .B2(KEYINPUT94), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(KEYINPUT94), .B2(new_n315_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n313_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n253_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n311_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n318_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n307_), .A2(new_n316_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n311_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n328_), .B1(new_n331_), .B2(new_n317_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n251_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n328_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n317_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n311_), .B1(new_n307_), .B2(new_n316_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n319_), .A2(new_n320_), .B1(new_n324_), .B2(new_n253_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n317_), .B(KEYINPUT27), .C1(new_n338_), .C2(new_n311_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(KEYINPUT96), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n333_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G141gat), .ZN(new_n344_));
  INV_X1    g143(.A(G148gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n343_), .A2(KEYINPUT2), .B1(new_n346_), .B2(KEYINPUT3), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n342_), .B(KEYINPUT82), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI221_X1 g148(.A(new_n347_), .B1(KEYINPUT3), .B2(new_n346_), .C1(new_n349_), .C2(KEYINPUT2), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  OR2_X1    g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(KEYINPUT1), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT83), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n352_), .B1(KEYINPUT1), .B2(new_n351_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n346_), .B(new_n348_), .C1(new_n355_), .C2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n295_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G78gat), .B(G106gat), .Z(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n364_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(KEYINPUT84), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n358_), .A2(new_n359_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT28), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n367_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n371_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G127gat), .B(G134gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G113gat), .B(G120gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n358_), .A2(KEYINPUT4), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n358_), .B(new_n378_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT4), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT92), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(KEYINPUT92), .A3(KEYINPUT4), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n375_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G85gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT0), .B(G57gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(new_n389_), .Z(new_n390_));
  INV_X1    g189(.A(new_n375_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n381_), .A2(new_n391_), .ZN(new_n392_));
  OR3_X1    g191(.A1(new_n386_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n390_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G15gat), .B(G43gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G71gat), .B(G99gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n303_), .B(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G227gat), .A2(G233gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n400_), .B(KEYINPUT80), .Z(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT30), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n399_), .B(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT81), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n403_), .A2(new_n404_), .ZN(new_n408_));
  MUX2_X1   g207(.A(new_n407_), .B(new_n406_), .S(new_n408_), .Z(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n395_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n341_), .A2(new_n374_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n395_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n372_), .A2(new_n373_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n337_), .A2(new_n413_), .A3(new_n414_), .A4(new_n339_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n381_), .A2(new_n391_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n417_), .A2(new_n390_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n384_), .A2(new_n375_), .A3(new_n385_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n384_), .A2(KEYINPUT93), .A3(new_n375_), .A4(new_n385_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n418_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n394_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n394_), .A2(new_n424_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n425_), .A2(new_n331_), .A3(new_n317_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n311_), .A2(KEYINPUT32), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n307_), .A2(new_n428_), .A3(new_n316_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n395_), .B(new_n429_), .C1(new_n338_), .C2(new_n428_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n414_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n410_), .B1(new_n416_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n250_), .B1(new_n412_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G230gat), .ZN(new_n434_));
  INV_X1    g233(.A(G233gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT66), .ZN(new_n437_));
  INV_X1    g236(.A(G57gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(G64gat), .ZN(new_n439_));
  INV_X1    g238(.A(G64gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(G57gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n437_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT11), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(G57gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n438_), .A2(G64gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(KEYINPUT66), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(new_n443_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT67), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G71gat), .B(G78gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n447_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n448_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n443_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n451_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n444_), .A2(new_n445_), .A3(KEYINPUT66), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT66), .B1(new_n444_), .B2(new_n445_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT11), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT67), .B1(new_n458_), .B2(new_n449_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n447_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n453_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n455_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G85gat), .B(G92gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT6), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(G99gat), .A3(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n464_), .B1(new_n468_), .B2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n463_), .B1(new_n474_), .B2(KEYINPUT65), .ZN(new_n475_));
  INV_X1    g274(.A(new_n464_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n470_), .A2(new_n472_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  INV_X1    g277(.A(G99gat), .ZN(new_n479_));
  INV_X1    g278(.A(G106gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n465_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n476_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n473_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n470_), .A2(new_n472_), .A3(KEYINPUT64), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n468_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n464_), .A2(KEYINPUT8), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n475_), .A2(new_n485_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT10), .B(G99gat), .Z(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n480_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n476_), .A2(KEYINPUT9), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n493_), .B(new_n494_), .C1(KEYINPUT9), .C2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n487_), .A2(new_n488_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n491_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n436_), .B1(new_n462_), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n454_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n459_), .A2(new_n460_), .A3(new_n453_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n489_), .A2(new_n490_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT8), .B1(new_n483_), .B2(new_n484_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n474_), .A2(KEYINPUT65), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n496_), .A2(new_n497_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT12), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n503_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n500_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n462_), .A2(new_n499_), .ZN(new_n515_));
  OAI22_X1  g314(.A1(new_n455_), .A2(new_n461_), .B1(new_n491_), .B2(new_n498_), .ZN(new_n516_));
  AOI211_X1 g315(.A(new_n434_), .B(new_n435_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G120gat), .B(G148gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G176gat), .B(G204gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n518_), .A2(new_n523_), .ZN(new_n526_));
  OR3_X1    g325(.A1(new_n525_), .A2(KEYINPUT13), .A3(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT13), .B1(new_n525_), .B2(new_n526_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G231gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n462_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(new_n227_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT76), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G127gat), .B(G155gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT16), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G183gat), .B(G211gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT17), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n533_), .B(new_n538_), .ZN(new_n539_));
  OR3_X1    g338(.A1(new_n532_), .A2(KEYINPUT17), .A3(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n499_), .A2(new_n206_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n509_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n543_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n547_), .A2(new_n548_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n551_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n543_), .A2(new_n544_), .A3(new_n553_), .A4(new_n549_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G190gat), .B(G218gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT70), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT72), .Z(new_n562_));
  NOR2_X1   g361(.A1(new_n555_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n555_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT73), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n559_), .B(KEYINPUT36), .Z(new_n566_));
  INV_X1    g365(.A(KEYINPUT73), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n555_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n563_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT37), .B1(new_n555_), .B2(new_n562_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n564_), .A2(new_n566_), .ZN(new_n571_));
  OAI22_X1  g370(.A1(new_n569_), .A2(KEYINPUT37), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n542_), .A2(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n433_), .A2(new_n529_), .A3(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(new_n207_), .A3(new_n395_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT38), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n569_), .B1(new_n412_), .B2(new_n432_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n529_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(new_n250_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n541_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT97), .Z(new_n582_));
  AND2_X1   g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(G1gat), .B1(new_n584_), .B2(new_n413_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n575_), .A2(new_n576_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n577_), .A2(new_n585_), .A3(new_n586_), .ZN(G1324gat));
  OAI21_X1  g386(.A(G8gat), .B1(new_n584_), .B2(new_n341_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT39), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n327_), .A2(new_n332_), .A3(new_n251_), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT96), .B1(new_n337_), .B2(new_n339_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n574_), .A2(new_n208_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT40), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(G1325gat));
  INV_X1    g395(.A(G15gat), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n574_), .A2(new_n597_), .A3(new_n409_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT98), .Z(new_n599_));
  AOI21_X1  g398(.A(new_n597_), .B1(new_n583_), .B2(new_n409_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT41), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n599_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(G1326gat));
  INV_X1    g405(.A(G22gat), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n583_), .B2(new_n414_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT42), .Z(new_n609_));
  NAND3_X1  g408(.A1(new_n574_), .A2(new_n607_), .A3(new_n414_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1327gat));
  NAND2_X1  g410(.A1(new_n580_), .A2(new_n542_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n411_), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n414_), .B(new_n613_), .C1(new_n333_), .C2(new_n340_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n431_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n409_), .B1(new_n615_), .B2(new_n415_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n572_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT43), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n572_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n572_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n412_), .B2(new_n432_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n612_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT44), .ZN(new_n627_));
  INV_X1    g426(.A(G29gat), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n413_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n630_));
  OAI211_X1 g429(.A(new_n627_), .B(new_n629_), .C1(new_n626_), .C2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n569_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n579_), .A2(new_n541_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n433_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n628_), .B1(new_n634_), .B2(new_n413_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n631_), .A2(new_n635_), .ZN(G1328gat));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT46), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n627_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G36gat), .B1(new_n641_), .B2(new_n341_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n341_), .A2(G36gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n433_), .A2(new_n633_), .A3(new_n643_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT102), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT102), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n645_), .A2(KEYINPUT45), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT45), .B1(new_n645_), .B2(new_n646_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n639_), .B(new_n640_), .C1(new_n642_), .C2(new_n649_), .ZN(new_n650_));
  AND4_X1   g449(.A1(new_n637_), .A2(new_n642_), .A3(new_n638_), .A4(new_n649_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1329gat));
  NAND2_X1  g451(.A1(new_n409_), .A2(G43gat), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n634_), .A2(new_n410_), .ZN(new_n654_));
  OAI22_X1  g453(.A1(new_n641_), .A2(new_n653_), .B1(G43gat), .B2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(G1330gat));
  NOR3_X1   g456(.A1(new_n634_), .A2(G50gat), .A3(new_n374_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n627_), .B(new_n414_), .C1(new_n626_), .C2(new_n630_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(G50gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT105), .ZN(G1331gat));
  NAND2_X1  g460(.A1(new_n579_), .A2(new_n250_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n542_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n578_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G57gat), .B1(new_n665_), .B2(new_n413_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n250_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT106), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT106), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n579_), .B(new_n573_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n395_), .A2(new_n438_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n670_), .B2(new_n671_), .ZN(G1332gat));
  AOI21_X1  g471(.A(new_n440_), .B1(new_n664_), .B2(new_n592_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT48), .Z(new_n674_));
  NAND2_X1  g473(.A1(new_n592_), .A2(new_n440_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n670_), .B2(new_n675_), .ZN(G1333gat));
  INV_X1    g475(.A(G71gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n664_), .B2(new_n409_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT107), .B(KEYINPUT49), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n409_), .A2(new_n677_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n670_), .B2(new_n681_), .ZN(G1334gat));
  INV_X1    g481(.A(G78gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n664_), .B2(new_n414_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n414_), .A2(new_n683_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n670_), .B2(new_n687_), .ZN(G1335gat));
  NOR2_X1   g487(.A1(new_n662_), .A2(new_n541_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G85gat), .B1(new_n692_), .B2(new_n413_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n541_), .A2(new_n632_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n579_), .B(new_n694_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n695_), .A2(new_n696_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n413_), .A2(G85gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n693_), .B1(new_n700_), .B2(new_n701_), .ZN(G1336gat));
  OAI21_X1  g501(.A(G92gat), .B1(new_n692_), .B2(new_n341_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n341_), .A2(G92gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n700_), .B2(new_n704_), .ZN(G1337gat));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(KEYINPUT111), .ZN(new_n707_));
  OAI21_X1  g506(.A(G99gat), .B1(new_n692_), .B2(new_n410_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT110), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n409_), .A2(new_n492_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n699_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n697_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n709_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n708_), .B(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n409_), .B(new_n492_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n707_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n713_), .A2(new_n718_), .ZN(G1338gat));
  OAI211_X1 g518(.A(new_n480_), .B(new_n414_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n623_), .A2(new_n624_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n622_), .B(new_n620_), .C1(new_n412_), .C2(new_n432_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n414_), .B(new_n689_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G106gat), .B1(new_n723_), .B2(KEYINPUT112), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n691_), .B2(new_n414_), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT52), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(KEYINPUT112), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n691_), .A2(new_n725_), .A3(new_n414_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n728_), .A2(new_n729_), .A3(new_n730_), .A4(G106gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n720_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT53), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n720_), .A2(new_n732_), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1339gat));
  INV_X1    g536(.A(KEYINPUT59), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n341_), .A2(new_n395_), .A3(new_n374_), .A4(new_n409_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n740_), .B2(KEYINPUT116), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(KEYINPUT116), .B2(new_n740_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n249_), .A2(new_n524_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT114), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n515_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n436_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n513_), .A2(KEYINPUT55), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n516_), .A2(KEYINPUT12), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n503_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n749_), .B1(new_n752_), .B2(new_n500_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n745_), .B(new_n747_), .C1(new_n748_), .C2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n523_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n513_), .A2(KEYINPUT55), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n752_), .A2(new_n749_), .A3(new_n500_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n745_), .B1(new_n760_), .B2(new_n747_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n756_), .A2(new_n757_), .A3(new_n761_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n758_), .A2(new_n759_), .B1(new_n436_), .B2(new_n746_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n523_), .B1(new_n763_), .B2(new_n745_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n747_), .B1(new_n748_), .B2(new_n753_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT114), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT56), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n744_), .B1(new_n762_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n243_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n233_), .A2(KEYINPUT78), .A3(new_n236_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n232_), .A2(new_n218_), .A3(new_n226_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n236_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n772_));
  AOI22_X1  g571(.A1(new_n769_), .A2(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n569_), .B1(new_n768_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT57), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n524_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n762_), .B2(new_n767_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT58), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n622_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n757_), .B1(new_n756_), .B2(new_n761_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n764_), .A2(KEYINPUT56), .A3(new_n766_), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n780_), .B(new_n777_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n743_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n774_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n632_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n781_), .A2(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n776_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n777_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n572_), .B1(new_n793_), .B2(KEYINPUT58), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n775_), .A2(KEYINPUT57), .B1(new_n794_), .B2(new_n784_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(KEYINPUT117), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n542_), .B1(new_n792_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT118), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n573_), .A2(new_n250_), .A3(new_n529_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n542_), .C1(new_n792_), .C2(new_n796_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n798_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n790_), .A2(new_n776_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n541_), .B1(new_n806_), .B2(KEYINPUT115), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(KEYINPUT115), .B2(new_n806_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n802_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n740_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n742_), .A2(new_n805_), .B1(new_n810_), .B2(KEYINPUT59), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n250_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n250_), .A2(G113gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n810_), .B2(new_n814_), .ZN(G1340gat));
  INV_X1    g614(.A(G120gat), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n811_), .B2(new_n579_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(KEYINPUT60), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n529_), .A2(KEYINPUT60), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n818_), .B(new_n810_), .C1(new_n816_), .C2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT119), .ZN(G1341gat));
  OAI21_X1  g621(.A(G127gat), .B1(new_n812_), .B2(new_n542_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n542_), .A2(G127gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n810_), .B2(new_n824_), .ZN(G1342gat));
  OAI21_X1  g624(.A(G134gat), .B1(new_n812_), .B2(new_n622_), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n632_), .A2(G134gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n810_), .B2(new_n827_), .ZN(G1343gat));
  AOI21_X1  g627(.A(new_n409_), .B1(new_n808_), .B2(new_n802_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(new_n395_), .A3(new_n414_), .A4(new_n341_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(new_n250_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(new_n344_), .ZN(G1344gat));
  NOR2_X1   g631(.A1(new_n830_), .A2(new_n529_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(new_n345_), .ZN(G1345gat));
  OR3_X1    g633(.A1(new_n830_), .A2(KEYINPUT120), .A3(new_n542_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT120), .B1(new_n830_), .B2(new_n542_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1346gat));
  OAI21_X1  g638(.A(G162gat), .B1(new_n830_), .B2(new_n622_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n632_), .A2(G162gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n830_), .B2(new_n841_), .ZN(G1347gat));
  NAND2_X1  g641(.A1(new_n592_), .A2(new_n411_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n414_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n795_), .A2(KEYINPUT117), .B1(KEYINPUT57), .B2(new_n775_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n790_), .A2(new_n791_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n541_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n802_), .B1(new_n847_), .B2(new_n803_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n804_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n844_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OR3_X1    g649(.A1(new_n850_), .A2(KEYINPUT121), .A3(new_n250_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT121), .B1(new_n850_), .B2(new_n250_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(G169gat), .A3(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT62), .ZN(new_n854_));
  INV_X1    g653(.A(new_n843_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n374_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n801_), .B1(new_n797_), .B2(KEYINPUT118), .ZN(new_n857_));
  AOI211_X1 g656(.A(KEYINPUT122), .B(new_n856_), .C1(new_n857_), .C2(new_n804_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n805_), .B2(new_n844_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n249_), .A2(new_n257_), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT123), .Z(new_n863_));
  OAI21_X1  g662(.A(new_n854_), .B1(new_n861_), .B2(new_n863_), .ZN(G1348gat));
  AOI21_X1  g663(.A(new_n414_), .B1(new_n808_), .B2(new_n802_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(G176gat), .A3(new_n579_), .A4(new_n855_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n850_), .A2(KEYINPUT122), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n805_), .A2(new_n859_), .A3(new_n844_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n529_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n258_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n869_), .A2(KEYINPUT124), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n579_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n258_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n866_), .B1(new_n871_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT125), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT125), .B(new_n866_), .C1(new_n871_), .C2(new_n874_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1349gat));
  NOR3_X1   g678(.A1(new_n861_), .A2(new_n268_), .A3(new_n542_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n843_), .A2(new_n542_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G183gat), .B1(new_n865_), .B2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n861_), .B2(new_n622_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n569_), .A2(new_n269_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n861_), .B2(new_n885_), .ZN(G1351gat));
  XNOR2_X1  g685(.A(KEYINPUT126), .B(G197gat), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(G197gat), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n341_), .A2(new_n395_), .A3(new_n374_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n829_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n250_), .ZN(new_n892_));
  MUX2_X1   g691(.A(new_n887_), .B(new_n889_), .S(new_n892_), .Z(G1352gat));
  INV_X1    g692(.A(new_n891_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n579_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n541_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  AND2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n897_), .B2(new_n898_), .ZN(G1354gat));
  AOI21_X1  g700(.A(G218gat), .B1(new_n894_), .B2(new_n569_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n572_), .A2(G218gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT127), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n894_), .B2(new_n904_), .ZN(G1355gat));
endmodule


