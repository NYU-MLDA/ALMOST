//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204_));
  AND2_X1   g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT7), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  AOI211_X1 g008(.A(new_n204_), .B(new_n205_), .C1(new_n207_), .C2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n203_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n213_), .B1(new_n210_), .B2(new_n203_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(KEYINPUT8), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT10), .B(G99gat), .Z(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(G92gat), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n204_), .B1(new_n205_), .B2(KEYINPUT9), .ZN(new_n227_));
  AND3_X1   g026(.A1(new_n226_), .A2(KEYINPUT66), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT66), .B1(new_n226_), .B2(new_n227_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n209_), .B(new_n220_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n217_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G29gat), .B(G36gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G43gat), .B(G50gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n230_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n230_), .A2(new_n236_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n237_), .A2(new_n238_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n234_), .B(KEYINPUT15), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n202_), .B(new_n235_), .C1(new_n239_), .C2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G232gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT73), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n239_), .A2(new_n241_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT35), .B1(new_n248_), .B2(new_n235_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n242_), .A2(new_n245_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n246_), .B(new_n247_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G190gat), .B(G218gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G134gat), .B(G162gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n254_), .A2(KEYINPUT36), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n251_), .B(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n249_), .A2(new_n250_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n246_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT36), .A3(new_n254_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT37), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT37), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n263_), .A3(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G15gat), .B(G22gat), .ZN(new_n266_));
  INV_X1    g065(.A(G1gat), .ZN(new_n267_));
  INV_X1    g066(.A(G8gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT14), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G1gat), .B(G8gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G231gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G57gat), .B(G64gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT11), .ZN(new_n276_));
  XOR2_X1   g075(.A(G71gat), .B(G78gat), .Z(new_n277_));
  OR2_X1    g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n275_), .A2(KEYINPUT11), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n277_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n274_), .B(new_n281_), .Z(new_n282_));
  XNOR2_X1  g081(.A(G127gat), .B(G155gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT16), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G183gat), .B(G211gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT17), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT74), .Z(new_n288_));
  NAND2_X1  g087(.A1(new_n282_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT75), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n286_), .B(KEYINPUT17), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n282_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n265_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT76), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G229gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n272_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n297_), .B1(new_n298_), .B2(new_n234_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n240_), .A2(new_n272_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n272_), .B(new_n234_), .Z(new_n301_));
  AOI22_X1  g100(.A1(new_n299_), .A2(new_n300_), .B1(new_n301_), .B2(new_n297_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G113gat), .B(G141gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G169gat), .B(G197gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT77), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n307_), .B(KEYINPUT78), .Z(new_n308_));
  NOR2_X1   g107(.A1(new_n302_), .A2(new_n305_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n231_), .A2(new_n281_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n231_), .A2(new_n281_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(KEYINPUT12), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n278_), .B(KEYINPUT12), .C1(new_n279_), .C2(new_n280_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n239_), .A2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(G230gat), .A2(G233gat), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n313_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n312_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n322_), .B(new_n317_), .C1(new_n321_), .C2(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G120gat), .B(G148gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT5), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G176gat), .B(G204gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n319_), .A2(new_n323_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT13), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(KEYINPUT71), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(KEYINPUT71), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n311_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G197gat), .A2(G204gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT89), .B(G204gat), .ZN(new_n339_));
  INV_X1    g138(.A(G197gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT21), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT91), .ZN(new_n343_));
  INV_X1    g142(.A(G211gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(G218gat), .ZN(new_n345_));
  INV_X1    g144(.A(G218gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(G211gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n343_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(G211gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(G218gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT91), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n341_), .A2(new_n342_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT90), .ZN(new_n353_));
  INV_X1    g152(.A(G204gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(G197gat), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(new_n339_), .B2(G197gat), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n354_), .A2(KEYINPUT89), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n354_), .A2(KEYINPUT89), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n353_), .B(new_n340_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(KEYINPUT21), .A3(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n348_), .A2(KEYINPUT21), .A3(new_n351_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n341_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n352_), .A2(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n368_));
  OR2_X1    g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(KEYINPUT3), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(KEYINPUT3), .B2(new_n369_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT87), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n367_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT88), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT88), .B(new_n367_), .C1(new_n371_), .C2(new_n373_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n366_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n365_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT86), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT85), .B1(new_n366_), .B2(KEYINPUT1), .ZN(new_n382_));
  OR3_X1    g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n383_), .B(new_n384_), .C1(KEYINPUT1), .C2(new_n366_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n386_));
  MUX2_X1   g185(.A(KEYINPUT84), .B(new_n386_), .S(new_n369_), .Z(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n378_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n363_), .B1(new_n389_), .B2(KEYINPUT29), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  XOR2_X1   g191(.A(G78gat), .B(G106gat), .Z(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT92), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT93), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n389_), .A2(KEYINPUT29), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G22gat), .B(G50gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT28), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n397_), .B(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n392_), .B(new_n394_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n401_), .A2(new_n402_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT27), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT18), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT23), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(G183gat), .B2(G190gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G183gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(KEYINPUT23), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT79), .B1(new_n417_), .B2(G190gat), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n413_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n415_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(KEYINPUT80), .A3(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT25), .B(G183gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT26), .B(G190gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G169gat), .A2(G176gat), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n425_), .A2(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n413_), .A2(G183gat), .A3(G190gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n414_), .B1(new_n434_), .B2(new_n419_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n431_), .B1(new_n435_), .B2(new_n422_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n424_), .A2(new_n430_), .A3(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT22), .B(G169gat), .ZN(new_n438_));
  INV_X1    g237(.A(G176gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n415_), .A2(new_n432_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n443_), .A2(new_n445_), .B1(G169gat), .B2(G176gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n363_), .A2(new_n437_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT95), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n421_), .A2(new_n449_), .A3(new_n445_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT95), .B1(new_n435_), .B2(new_n444_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n429_), .B(KEYINPUT94), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n439_), .B2(new_n438_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n430_), .A2(new_n443_), .A3(new_n423_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(KEYINPUT20), .B(new_n448_), .C1(new_n456_), .C2(new_n363_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT96), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G226gat), .A2(G233gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT19), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n363_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n460_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n437_), .A2(new_n447_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n363_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n462_), .A2(KEYINPUT20), .A3(new_n463_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n461_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n458_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n469_));
  OAI211_X1 g268(.A(KEYINPUT98), .B(new_n412_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n363_), .A2(new_n437_), .A3(new_n447_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n352_), .A2(new_n360_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n361_), .A2(new_n362_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n454_), .A2(new_n455_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n472_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT96), .B1(new_n477_), .B2(new_n463_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n467_), .A3(new_n461_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT98), .B1(new_n479_), .B2(new_n412_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n471_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n468_), .A2(new_n469_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(KEYINPUT97), .A3(new_n411_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n478_), .A2(new_n411_), .A3(new_n467_), .A4(new_n461_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT97), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n407_), .B1(new_n481_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n462_), .A2(KEYINPUT20), .A3(new_n466_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n460_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n460_), .B2(new_n457_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n412_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(KEYINPUT27), .A3(new_n484_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n406_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G127gat), .B(G134gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G113gat), .B(G120gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n378_), .A2(new_n388_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n378_), .B2(new_n388_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G225gat), .A2(G233gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n500_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n389_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n378_), .A2(new_n388_), .A3(new_n500_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(KEYINPUT4), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n502_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n507_), .B1(new_n514_), .B2(new_n504_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G1gat), .B(G29gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(G85gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT0), .B(G57gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  OR2_X1    g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n519_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G227gat), .A2(G233gat), .ZN(new_n524_));
  INV_X1    g323(.A(G71gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G99gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n464_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n500_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G15gat), .B(G43gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT82), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT30), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT31), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n529_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n495_), .A2(new_n523_), .A3(new_n536_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n405_), .A2(new_n522_), .A3(new_n494_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n491_), .A2(KEYINPUT32), .A3(new_n411_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n411_), .A2(KEYINPUT32), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n482_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT101), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n540_), .A2(new_n543_), .A3(KEYINPUT102), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT102), .B1(new_n540_), .B2(new_n543_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT99), .B1(new_n481_), .B2(new_n487_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n412_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT98), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n470_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT99), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(new_n486_), .A4(new_n483_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n514_), .A2(new_n504_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n519_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n503_), .A2(new_n505_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT33), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n515_), .B2(new_n519_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n504_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n559_), .B(new_n519_), .C1(new_n561_), .C2(new_n506_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n558_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT100), .B1(new_n554_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT100), .ZN(new_n567_));
  AOI211_X1 g366(.A(new_n567_), .B(new_n564_), .C1(new_n547_), .C2(new_n553_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n546_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n538_), .B1(new_n569_), .B2(new_n405_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n537_), .B1(new_n570_), .B2(new_n536_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n336_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n295_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n267_), .A3(new_n522_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT38), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n571_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n261_), .B(KEYINPUT103), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n293_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n336_), .A3(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G1gat), .B1(new_n582_), .B2(new_n523_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n574_), .A2(new_n575_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n576_), .A2(new_n583_), .A3(new_n584_), .ZN(G1324gat));
  NAND3_X1  g384(.A1(new_n573_), .A2(new_n268_), .A3(new_n494_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n494_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n582_), .A2(KEYINPUT104), .A3(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(new_n268_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT104), .B1(new_n582_), .B2(new_n587_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n586_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT40), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(KEYINPUT40), .B(new_n586_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(G1325gat));
  INV_X1    g397(.A(new_n536_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G15gat), .B1(new_n582_), .B2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT41), .Z(new_n601_));
  INV_X1    g400(.A(G15gat), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n573_), .A2(new_n602_), .A3(new_n536_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT105), .ZN(G1326gat));
  OAI21_X1  g404(.A(G22gat), .B1(new_n582_), .B2(new_n405_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT42), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n405_), .A2(G22gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT106), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n573_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(G1327gat));
  INV_X1    g410(.A(new_n261_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(new_n581_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n572_), .A2(new_n613_), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n614_), .A2(G29gat), .A3(new_n523_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT43), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n569_), .A2(new_n405_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n538_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n536_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n537_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n616_), .B(new_n265_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT107), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT107), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n571_), .A2(new_n623_), .A3(new_n616_), .A4(new_n265_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n571_), .A2(new_n265_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT43), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n622_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n336_), .A2(new_n293_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT44), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n627_), .A2(new_n628_), .A3(KEYINPUT44), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n631_), .A2(KEYINPUT108), .A3(new_n522_), .A4(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(G29gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n631_), .A2(new_n522_), .A3(new_n632_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT108), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT109), .B1(new_n634_), .B2(new_n637_), .ZN(new_n638_));
  AND4_X1   g437(.A1(KEYINPUT109), .A2(new_n637_), .A3(G29gat), .A4(new_n633_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n615_), .B1(new_n638_), .B2(new_n639_), .ZN(G1328gat));
  NOR2_X1   g439(.A1(new_n587_), .A2(G36gat), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n336_), .A2(new_n571_), .A3(new_n613_), .A4(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n642_), .B(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n631_), .A2(new_n494_), .A3(new_n632_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(G36gat), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT111), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n648_), .B(new_n651_), .ZN(G1329gat));
  AND3_X1   g451(.A1(new_n631_), .A2(new_n536_), .A3(new_n632_), .ZN(new_n653_));
  INV_X1    g452(.A(G43gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n536_), .A2(new_n654_), .ZN(new_n655_));
  OAI22_X1  g454(.A1(new_n653_), .A2(new_n654_), .B1(new_n614_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT47), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(G1330gat));
  OR3_X1    g457(.A1(new_n614_), .A2(G50gat), .A3(new_n405_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n631_), .A2(new_n406_), .A3(new_n632_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(KEYINPUT112), .A3(G50gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT112), .B1(new_n660_), .B2(G50gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(G1331gat));
  NAND2_X1  g462(.A1(new_n334_), .A2(new_n335_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(new_n310_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(new_n293_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(new_n580_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G57gat), .B1(new_n669_), .B2(new_n523_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n666_), .A2(new_n577_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(new_n295_), .ZN(new_n672_));
  INV_X1    g471(.A(G57gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n522_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n674_), .ZN(G1332gat));
  INV_X1    g474(.A(G64gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n672_), .A2(new_n676_), .A3(new_n494_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n668_), .A2(new_n494_), .ZN(new_n678_));
  XOR2_X1   g477(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n679_));
  AND3_X1   g478(.A1(new_n678_), .A2(G64gat), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n678_), .B2(G64gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(G1333gat));
  AOI21_X1  g481(.A(new_n525_), .B1(new_n668_), .B2(new_n536_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT49), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n672_), .A2(new_n525_), .A3(new_n536_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1334gat));
  INV_X1    g485(.A(G78gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n668_), .B2(new_n406_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT50), .Z(new_n689_));
  NAND3_X1  g488(.A1(new_n672_), .A2(new_n687_), .A3(new_n406_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1335gat));
  AND3_X1   g490(.A1(new_n627_), .A2(new_n293_), .A3(new_n665_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G85gat), .B1(new_n693_), .B2(new_n523_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n671_), .A2(new_n613_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n223_), .A3(new_n522_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1336gat));
  AOI21_X1  g496(.A(G92gat), .B1(new_n695_), .B2(new_n494_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n587_), .A2(new_n222_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n692_), .B2(new_n699_), .ZN(G1337gat));
  NAND2_X1  g499(.A1(new_n692_), .A2(new_n536_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n536_), .A2(new_n218_), .ZN(new_n702_));
  AOI22_X1  g501(.A1(new_n701_), .A2(G99gat), .B1(new_n695_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g503(.A1(new_n695_), .A2(new_n219_), .A3(new_n406_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n627_), .A2(new_n293_), .A3(new_n406_), .A4(new_n665_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G106gat), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT52), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(KEYINPUT52), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n705_), .B(new_n706_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n708_), .B(KEYINPUT52), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n706_), .B1(new_n713_), .B2(new_n705_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1339gat));
  NAND3_X1  g514(.A1(new_n294_), .A2(new_n311_), .A3(new_n333_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT54), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n310_), .A2(new_n331_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT55), .B1(new_n318_), .B2(KEYINPUT115), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT115), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT55), .ZN(new_n722_));
  OAI221_X1 g521(.A(new_n312_), .B1(new_n313_), .B2(KEYINPUT12), .C1(new_n239_), .C2(new_n315_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n721_), .B(new_n722_), .C1(new_n723_), .C2(new_n317_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n317_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n720_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT56), .B1(new_n726_), .B2(new_n328_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n726_), .A2(KEYINPUT56), .A3(new_n328_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n719_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n305_), .B1(new_n301_), .B2(new_n296_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n732_), .A2(KEYINPUT116), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n296_), .B1(new_n298_), .B2(new_n234_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n732_), .A2(KEYINPUT116), .B1(new_n300_), .B2(new_n734_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n733_), .A2(new_n735_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n332_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n612_), .B1(new_n730_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT57), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT117), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n729_), .A2(new_n741_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n726_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n328_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n728_), .A3(new_n743_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n331_), .A2(new_n736_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(KEYINPUT58), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n265_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT58), .B1(new_n744_), .B2(new_n745_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n581_), .B1(new_n740_), .B2(new_n749_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n718_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT120), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(KEYINPUT59), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n495_), .A2(new_n522_), .A3(new_n536_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT119), .ZN(new_n755_));
  MUX2_X1   g554(.A(new_n752_), .B(new_n753_), .S(new_n755_), .Z(new_n756_));
  NAND2_X1  g555(.A1(new_n751_), .A2(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n739_), .A2(KEYINPUT57), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n739_), .A2(KEYINPUT57), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n758_), .A2(new_n759_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT118), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT118), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n740_), .A2(new_n749_), .A3(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n761_), .A2(new_n293_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n718_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(new_n755_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT59), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n757_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G113gat), .B1(new_n769_), .B2(new_n311_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n766_), .A2(new_n755_), .ZN(new_n771_));
  OR3_X1    g570(.A1(new_n771_), .A2(G113gat), .A3(new_n311_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1340gat));
  OAI21_X1  g572(.A(G120gat), .B1(new_n769_), .B2(new_n664_), .ZN(new_n774_));
  INV_X1    g573(.A(G120gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n664_), .B2(KEYINPUT60), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n767_), .B(new_n776_), .C1(KEYINPUT60), .C2(new_n775_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(G1341gat));
  OAI21_X1  g577(.A(G127gat), .B1(new_n769_), .B2(new_n293_), .ZN(new_n779_));
  OR3_X1    g578(.A1(new_n771_), .A2(G127gat), .A3(new_n293_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1342gat));
  AOI21_X1  g580(.A(G134gat), .B1(new_n767_), .B2(new_n579_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n769_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n265_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT121), .B(G134gat), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n782_), .B1(new_n783_), .B2(new_n786_), .ZN(G1343gat));
  NOR2_X1   g586(.A1(new_n405_), .A2(new_n536_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n494_), .A2(new_n523_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n766_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n310_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g591(.A(new_n664_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g594(.A(KEYINPUT61), .B(G155gat), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n766_), .A2(new_n581_), .A3(new_n788_), .A4(new_n789_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(KEYINPUT122), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(KEYINPUT122), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n797_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n798_), .A2(KEYINPUT122), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n798_), .A2(KEYINPUT122), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n796_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(G1346gat));
  INV_X1    g604(.A(new_n790_), .ZN(new_n806_));
  OAI21_X1  g605(.A(G162gat), .B1(new_n806_), .B2(new_n784_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n578_), .A2(G162gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n806_), .B2(new_n808_), .ZN(G1347gat));
  NOR2_X1   g608(.A1(new_n587_), .A2(new_n522_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(new_n599_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n311_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n751_), .A2(new_n405_), .A3(new_n438_), .A4(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT123), .B1(new_n813_), .B2(new_n311_), .ZN(new_n816_));
  OR3_X1    g615(.A1(new_n813_), .A2(KEYINPUT123), .A3(new_n311_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n751_), .A2(new_n405_), .A3(new_n816_), .A4(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(G169gat), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n818_), .B2(G169gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n815_), .B1(new_n821_), .B2(new_n822_), .ZN(G1348gat));
  NAND3_X1  g622(.A1(new_n751_), .A2(new_n405_), .A3(new_n812_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n439_), .B1(new_n824_), .B2(new_n664_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n406_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n826_), .A2(G176gat), .A3(new_n793_), .A4(new_n812_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT124), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n825_), .A2(new_n830_), .A3(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1349gat));
  NOR3_X1   g631(.A1(new_n824_), .A2(new_n293_), .A3(new_n425_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n826_), .A2(new_n581_), .A3(new_n812_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n416_), .B2(new_n834_), .ZN(G1350gat));
  OAI21_X1  g634(.A(G190gat), .B1(new_n824_), .B2(new_n784_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n579_), .A2(new_n426_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n824_), .B2(new_n837_), .ZN(G1351gat));
  AND3_X1   g637(.A1(new_n766_), .A2(new_n788_), .A3(new_n810_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n310_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g640(.A1(new_n766_), .A2(new_n793_), .A3(new_n788_), .A4(new_n810_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n843_));
  INV_X1    g642(.A(new_n339_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n842_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n842_), .A2(new_n844_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(KEYINPUT125), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n842_), .A2(G204gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n845_), .B1(new_n847_), .B2(new_n848_), .ZN(G1353gat));
  AOI21_X1  g648(.A(new_n293_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT126), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n839_), .A2(new_n851_), .ZN(new_n852_));
  OR2_X1    g651(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1354gat));
  AOI21_X1  g653(.A(G218gat), .B1(new_n839_), .B2(new_n579_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n265_), .A2(G218gat), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT127), .Z(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n839_), .B2(new_n857_), .ZN(G1355gat));
endmodule


