//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_;
  NOR2_X1   g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  AND3_X1   g004(.A1(new_n205_), .A2(KEYINPUT64), .A3(new_n204_), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT64), .B1(new_n205_), .B2(new_n204_), .ZN(new_n207_));
  OAI221_X1 g006(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .C1(new_n206_), .C2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT6), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT10), .B(G99gat), .Z(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(new_n210_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n208_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n211_), .A2(KEYINPUT65), .A3(new_n213_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT65), .B1(new_n211_), .B2(new_n213_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT66), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n221_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n219_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT7), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n203_), .A2(new_n205_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n218_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  AOI211_X1 g030(.A(KEYINPUT8), .B(new_n229_), .C1(new_n227_), .C2(new_n214_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n217_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G29gat), .B(G36gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G43gat), .B(G50gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT15), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n236_), .B(new_n217_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G232gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT34), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT35), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n238_), .A2(new_n239_), .A3(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n242_), .A2(new_n243_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n245_), .A2(new_n246_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G190gat), .B(G218gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G134gat), .B(G162gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  OR4_X1    g050(.A1(KEYINPUT36), .A2(new_n247_), .A3(new_n248_), .A4(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(KEYINPUT36), .Z(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(KEYINPUT37), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT37), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G57gat), .B(G64gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT11), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n260_), .A2(KEYINPUT11), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT67), .B(G71gat), .ZN(new_n265_));
  INV_X1    g064(.A(G78gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n261_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G15gat), .B(G22gat), .ZN(new_n271_));
  INV_X1    g070(.A(G1gat), .ZN(new_n272_));
  INV_X1    g071(.A(G8gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT14), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G1gat), .B(G8gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G231gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n270_), .B(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G127gat), .B(G155gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(G183gat), .B(G211gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT70), .B(KEYINPUT16), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT17), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(KEYINPUT17), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n280_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT72), .Z(new_n289_));
  NOR2_X1   g088(.A1(new_n280_), .A2(new_n286_), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n290_), .B(KEYINPUT71), .Z(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n259_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT73), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n270_), .B(new_n217_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n270_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n233_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(G230gat), .A2(G233gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n296_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(new_n302_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT12), .B1(new_n300_), .B2(KEYINPUT69), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT69), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT12), .ZN(new_n308_));
  AOI211_X1 g107(.A(new_n307_), .B(new_n308_), .C1(new_n233_), .C2(new_n299_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n305_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n303_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G120gat), .B(G148gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT5), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G176gat), .B(G204gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n303_), .A2(new_n310_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT13), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT13), .B1(new_n316_), .B2(new_n318_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n295_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G134gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G127gat), .ZN(new_n327_));
  INV_X1    g126(.A(G127gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G134gat), .ZN(new_n329_));
  INV_X1    g128(.A(G120gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(G113gat), .ZN(new_n331_));
  INV_X1    g130(.A(G113gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G120gat), .ZN(new_n333_));
  AND4_X1   g132(.A1(new_n327_), .A2(new_n329_), .A3(new_n331_), .A4(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n327_), .A2(new_n329_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT31), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(KEYINPUT23), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(KEYINPUT23), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n343_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G183gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT25), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G183gat), .ZN(new_n355_));
  INV_X1    g154(.A(G190gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT26), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT26), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(G190gat), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n353_), .A2(new_n355_), .A3(new_n357_), .A4(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n347_), .B1(G169gat), .B2(G176gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n346_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT78), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n345_), .A2(KEYINPUT80), .A3(new_n348_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n360_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n351_), .A2(new_n365_), .A3(new_n366_), .A4(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n343_), .A2(G183gat), .A3(G190gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n342_), .A2(new_n370_), .A3(KEYINPUT81), .ZN(new_n371_));
  OR3_X1    g170(.A1(new_n340_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n352_), .A2(new_n356_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n371_), .A2(new_n372_), .A3(KEYINPUT82), .A4(new_n373_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G169gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n369_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382_));
  INV_X1    g181(.A(G71gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G99gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n381_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G15gat), .B(G43gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT83), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n388_), .B(KEYINPUT30), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n386_), .B(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n338_), .B1(new_n390_), .B2(KEYINPUT84), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(KEYINPUT84), .B2(new_n390_), .ZN(new_n392_));
  OR3_X1    g191(.A1(new_n390_), .A2(KEYINPUT84), .A3(new_n337_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n399_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G141gat), .ZN(new_n409_));
  INV_X1    g208(.A(G148gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n396_), .B1(KEYINPUT1), .B2(new_n398_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT1), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(G155gat), .A3(G162gat), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n413_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n336_), .B1(new_n408_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT2), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n412_), .A2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n420_), .A2(new_n422_), .A3(new_n404_), .A4(new_n400_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n398_), .A3(new_n397_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n327_), .A2(new_n329_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n331_), .A2(new_n333_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n327_), .A2(new_n329_), .A3(new_n331_), .A4(new_n333_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n398_), .A2(KEYINPUT1), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n397_), .A2(new_n430_), .A3(new_n416_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n424_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n418_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n435_), .B(KEYINPUT90), .Z(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n418_), .A2(KEYINPUT4), .A3(new_n433_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n418_), .A2(new_n433_), .A3(KEYINPUT89), .A4(KEYINPUT4), .ZN(new_n441_));
  INV_X1    g240(.A(new_n418_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n437_), .B1(new_n445_), .B2(new_n436_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G57gat), .B(G85gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n446_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n451_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n436_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n438_), .A2(new_n439_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n455_), .B2(new_n441_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n453_), .B1(new_n456_), .B2(new_n437_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n458_), .A2(KEYINPUT95), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(KEYINPUT95), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n395_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT97), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G226gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT19), .ZN(new_n466_));
  OR2_X1    g265(.A1(G197gat), .A2(G204gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G197gat), .A2(G204gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G211gat), .B(G218gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n470_), .A2(new_n472_), .A3(KEYINPUT86), .A4(KEYINPUT21), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT86), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n467_), .A2(KEYINPUT21), .A3(new_n468_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n474_), .B1(new_n475_), .B2(new_n471_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n475_), .A2(new_n471_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT21), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n469_), .A2(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n473_), .A2(new_n476_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n369_), .A2(new_n380_), .A3(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n361_), .A2(KEYINPUT88), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n361_), .A2(KEYINPUT88), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n362_), .A3(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n371_), .A2(new_n372_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n348_), .A4(new_n360_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n345_), .A2(new_n373_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n379_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n480_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n482_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT87), .B1(new_n481_), .B2(KEYINPUT20), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n466_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n487_), .A2(new_n480_), .A3(new_n489_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT20), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n480_), .B1(new_n369_), .B2(new_n380_), .ZN(new_n498_));
  OR3_X1    g297(.A1(new_n497_), .A2(new_n498_), .A3(new_n466_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G8gat), .B(G36gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT18), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G64gat), .B(G92gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT27), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n495_), .A2(new_n504_), .A3(new_n499_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(KEYINPUT96), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT93), .B(new_n466_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n466_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n481_), .A2(KEYINPUT20), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(new_n492_), .A3(new_n482_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n512_), .B(new_n515_), .C1(new_n519_), .C2(new_n466_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n505_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT96), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n495_), .A2(new_n522_), .A3(new_n504_), .A4(new_n499_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n511_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n510_), .B1(KEYINPUT27), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n424_), .A2(new_n432_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT29), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n491_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G22gat), .B(G50gat), .Z(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n526_), .A2(KEYINPUT29), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n532_), .A2(KEYINPUT28), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT85), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(KEYINPUT28), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G228gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(new_n266_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n210_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n534_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n537_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n540_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n532_), .B(KEYINPUT28), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT85), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n545_), .B2(new_n536_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n531_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n540_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n543_), .A3(new_n536_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n530_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n464_), .B1(new_n525_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n524_), .A2(KEYINPUT27), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n509_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n551_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(KEYINPUT97), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n463_), .B1(new_n552_), .B2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT33), .B1(new_n446_), .B2(new_n451_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT33), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n559_), .B(new_n453_), .C1(new_n456_), .C2(new_n437_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n455_), .A2(new_n454_), .A3(new_n441_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n453_), .B1(new_n436_), .B2(new_n434_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n506_), .A2(new_n561_), .A3(new_n508_), .A4(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n558_), .A2(new_n560_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n568_), .A2(KEYINPUT92), .A3(new_n508_), .A4(new_n506_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n504_), .A2(KEYINPUT32), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n520_), .A2(new_n570_), .B1(new_n457_), .B2(new_n452_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n500_), .A2(new_n570_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n567_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n555_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT94), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n565_), .A2(new_n566_), .B1(new_n572_), .B2(new_n571_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n551_), .B1(new_n577_), .B2(new_n569_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n554_), .A2(new_n551_), .A3(new_n462_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n576_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n557_), .B1(new_n582_), .B2(new_n394_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G113gat), .B(G141gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT77), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G169gat), .B(G197gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n585_), .B(new_n586_), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n236_), .B(KEYINPUT74), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(new_n277_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT75), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n237_), .A2(new_n277_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT76), .ZN(new_n595_));
  INV_X1    g394(.A(new_n277_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n592_), .B1(new_n588_), .B2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n587_), .B1(new_n593_), .B2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n587_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n583_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n325_), .A2(new_n605_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n606_), .A2(G1gat), .A3(new_n462_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n608_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n255_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n583_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n323_), .A2(new_n603_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n292_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n461_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G1gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n609_), .A2(new_n610_), .A3(new_n616_), .ZN(G1324gat));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n525_), .A3(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(G8gat), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(KEYINPUT39), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(KEYINPUT39), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n525_), .A2(new_n273_), .ZN(new_n622_));
  OAI22_X1  g421(.A1(new_n620_), .A2(new_n621_), .B1(new_n606_), .B2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g423(.A1(new_n606_), .A2(G15gat), .A3(new_n394_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n612_), .A2(new_n395_), .A3(new_n614_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n626_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT41), .B1(new_n626_), .B2(G15gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT99), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n625_), .B(new_n631_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(G1326gat));
  OR3_X1    g432(.A1(new_n606_), .A2(G22gat), .A3(new_n555_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n612_), .A2(new_n551_), .A3(new_n614_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(G22gat), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(KEYINPUT42), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n636_), .A2(KEYINPUT42), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n634_), .B(KEYINPUT100), .C1(new_n638_), .C2(new_n637_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1327gat));
  NAND2_X1  g442(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n551_), .B1(new_n460_), .B2(new_n459_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n509_), .B2(new_n553_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n575_), .B2(KEYINPUT94), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n395_), .B1(new_n647_), .B2(new_n580_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n644_), .B1(new_n648_), .B2(new_n557_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n256_), .A2(new_n258_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n581_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n575_), .A2(KEYINPUT94), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n394_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n557_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(KEYINPUT102), .A3(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n649_), .A2(new_n650_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(KEYINPUT101), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n657_), .A2(KEYINPUT101), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n583_), .B2(new_n259_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n613_), .A2(new_n293_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n656_), .A2(new_n659_), .A3(new_n661_), .A4(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n650_), .B1(new_n648_), .B2(new_n557_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n658_), .B1(new_n666_), .B2(new_n660_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(new_n656_), .A3(KEYINPUT44), .A4(new_n662_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n665_), .A2(new_n668_), .A3(G29gat), .A4(new_n461_), .ZN(new_n669_));
  INV_X1    g468(.A(G29gat), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n255_), .A2(new_n293_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n324_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n605_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n674_), .B2(new_n462_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n669_), .A2(new_n675_), .ZN(G1328gat));
  NAND3_X1  g475(.A1(new_n665_), .A2(new_n525_), .A3(new_n668_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n554_), .A2(G36gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n679_), .B1(new_n674_), .B2(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n605_), .A2(KEYINPUT45), .A3(new_n673_), .A4(new_n680_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n678_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n687_));
  NOR2_X1   g486(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT104), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n686_), .A2(new_n687_), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n689_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n684_), .B1(new_n677_), .B2(G36gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n687_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(new_n694_), .ZN(G1329gat));
  NAND4_X1  g494(.A1(new_n665_), .A2(new_n668_), .A3(G43gat), .A4(new_n395_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n674_), .A2(new_n394_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(G43gat), .B2(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(G1330gat));
  NAND4_X1  g499(.A1(new_n665_), .A2(new_n668_), .A3(G50gat), .A4(new_n551_), .ZN(new_n701_));
  INV_X1    g500(.A(G50gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n674_), .B2(new_n555_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1331gat));
  NOR3_X1   g503(.A1(new_n323_), .A2(new_n603_), .A3(new_n292_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT107), .B(G57gat), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n612_), .A2(new_n461_), .A3(new_n705_), .A4(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT108), .Z(new_n708_));
  NOR2_X1   g507(.A1(new_n295_), .A2(new_n323_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n583_), .A2(new_n603_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n462_), .B1(new_n711_), .B2(KEYINPUT106), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(KEYINPUT106), .B2(new_n711_), .ZN(new_n713_));
  INV_X1    g512(.A(G57gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n708_), .B1(new_n713_), .B2(new_n714_), .ZN(G1332gat));
  NAND3_X1  g514(.A1(new_n612_), .A2(new_n525_), .A3(new_n705_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(G64gat), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(G64gat), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n554_), .A2(G64gat), .ZN(new_n720_));
  OAI22_X1  g519(.A1(new_n718_), .A2(new_n719_), .B1(new_n711_), .B2(new_n720_), .ZN(G1333gat));
  NAND3_X1  g520(.A1(new_n612_), .A2(new_n395_), .A3(new_n705_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G71gat), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT49), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n395_), .A2(new_n383_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n711_), .B2(new_n725_), .ZN(G1334gat));
  NAND3_X1  g525(.A1(new_n612_), .A2(new_n551_), .A3(new_n705_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(G78gat), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G78gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n551_), .A2(new_n266_), .ZN(new_n731_));
  OAI22_X1  g530(.A1(new_n729_), .A2(new_n730_), .B1(new_n711_), .B2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT111), .Z(G1335gat));
  NAND2_X1  g532(.A1(new_n667_), .A2(new_n656_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n604_), .A2(new_n292_), .ZN(new_n737_));
  OR3_X1    g536(.A1(new_n323_), .A2(KEYINPUT113), .A3(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT113), .B1(new_n323_), .B2(new_n737_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n736_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n667_), .A2(KEYINPUT112), .A3(new_n656_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n461_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G85gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n323_), .A2(new_n672_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n710_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n462_), .A2(G85gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1336gat));
  NAND3_X1  g548(.A1(new_n741_), .A2(new_n525_), .A3(new_n742_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G92gat), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n554_), .A2(G92gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n747_), .B2(new_n752_), .ZN(G1337gat));
  NAND4_X1  g552(.A1(new_n736_), .A2(new_n395_), .A3(new_n742_), .A4(new_n740_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G99gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n746_), .A2(new_n395_), .A3(new_n215_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT51), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n759_), .A3(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1338gat));
  AOI21_X1  g560(.A(new_n555_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n656_), .A2(new_n762_), .A3(new_n659_), .A4(new_n661_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n667_), .A2(new_n656_), .A3(KEYINPUT114), .A4(new_n762_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(G106gat), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(KEYINPUT52), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n765_), .A2(new_n766_), .A3(G106gat), .A4(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n746_), .A2(new_n210_), .A3(new_n551_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT53), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n770_), .A2(new_n776_), .A3(new_n772_), .A4(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1339gat));
  NAND4_X1  g577(.A1(new_n259_), .A2(new_n604_), .A3(new_n323_), .A4(new_n293_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT54), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n298_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n302_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n310_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT55), .B(new_n305_), .C1(new_n306_), .C2(new_n309_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n787_));
  OR2_X1    g586(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n786_), .A2(new_n315_), .A3(new_n787_), .A4(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n590_), .A2(new_n591_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n591_), .B1(new_n588_), .B2(new_n596_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n601_), .B1(new_n595_), .B2(new_n791_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n600_), .A2(new_n601_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n318_), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n302_), .A2(new_n781_), .B1(new_n310_), .B2(new_n783_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n317_), .B1(new_n795_), .B2(new_n785_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n789_), .B(new_n794_), .C1(new_n796_), .C2(new_n787_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n786_), .A2(new_n315_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n801_), .A2(KEYINPUT58), .A3(new_n789_), .A4(new_n794_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n650_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n796_), .B2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n800_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n603_), .A2(new_n318_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n807_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n319_), .A2(new_n793_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n611_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n803_), .B1(new_n812_), .B2(KEYINPUT57), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n814_), .B(new_n611_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n292_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n780_), .A2(new_n816_), .ZN(new_n817_));
  AOI211_X1 g616(.A(new_n394_), .B(new_n462_), .C1(new_n552_), .C2(new_n556_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n332_), .B1(new_n819_), .B2(new_n604_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT118), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n820_), .A2(KEYINPUT118), .ZN(new_n822_));
  INV_X1    g621(.A(new_n819_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  INV_X1    g623(.A(new_n780_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n816_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT119), .B(new_n292_), .C1(new_n813_), .C2(new_n815_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n825_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n818_), .A2(new_n824_), .ZN(new_n830_));
  OAI22_X1  g629(.A1(new_n823_), .A2(new_n824_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n603_), .A2(G113gat), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT120), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n821_), .A2(new_n822_), .B1(new_n832_), .B2(new_n834_), .ZN(G1340gat));
  XOR2_X1   g634(.A(KEYINPUT121), .B(G120gat), .Z(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n831_), .B2(new_n323_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n323_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(KEYINPUT60), .B2(new_n836_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n819_), .B2(new_n840_), .ZN(G1341gat));
  AOI21_X1  g640(.A(G127gat), .B1(new_n823_), .B2(new_n293_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n328_), .B1(new_n293_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n843_), .B2(new_n328_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n832_), .B2(new_n845_), .ZN(G1342gat));
  OAI21_X1  g645(.A(G134gat), .B1(new_n831_), .B2(new_n259_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n823_), .A2(new_n326_), .A3(new_n611_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1343gat));
  AOI21_X1  g648(.A(new_n395_), .B1(new_n780_), .B2(new_n816_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(new_n551_), .A3(new_n461_), .A4(new_n554_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n604_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(new_n409_), .ZN(G1344gat));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n323_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT123), .B(G148gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1345gat));
  NOR2_X1   g655(.A1(new_n851_), .A2(new_n292_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT61), .B(G155gat), .Z(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1346gat));
  OAI21_X1  g658(.A(G162gat), .B1(new_n851_), .B2(new_n259_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n255_), .A2(G162gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n851_), .B2(new_n861_), .ZN(G1347gat));
  NAND2_X1  g661(.A1(new_n800_), .A2(KEYINPUT116), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n808_), .B1(new_n863_), .B2(new_n804_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n864_), .A2(new_n807_), .B1(new_n319_), .B2(new_n793_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n814_), .B1(new_n865_), .B2(new_n611_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n812_), .A2(KEYINPUT57), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n803_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT119), .B1(new_n868_), .B2(new_n292_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n828_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n780_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT22), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n463_), .A2(new_n554_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n551_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n871_), .A2(new_n872_), .A3(new_n603_), .A4(new_n875_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(G169gat), .A3(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n876_), .A2(new_n878_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n871_), .A2(new_n603_), .A3(new_n877_), .A4(new_n875_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(G169gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n879_), .B1(new_n880_), .B2(new_n882_), .ZN(G1348gat));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884_));
  INV_X1    g683(.A(new_n875_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n827_), .A2(new_n828_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n780_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G176gat), .B1(new_n887_), .B2(new_n324_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n324_), .A2(G176gat), .A3(new_n873_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n817_), .A2(new_n555_), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n884_), .B1(new_n888_), .B2(new_n891_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n829_), .A2(new_n323_), .A3(new_n885_), .ZN(new_n893_));
  OAI211_X1 g692(.A(KEYINPUT125), .B(new_n890_), .C1(new_n893_), .C2(G176gat), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1349gat));
  AND4_X1   g694(.A1(new_n555_), .A2(new_n817_), .A3(new_n293_), .A4(new_n873_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(G183gat), .B1(new_n896_), .B2(new_n897_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n292_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n898_), .A2(new_n899_), .B1(new_n887_), .B2(new_n900_), .ZN(G1350gat));
  INV_X1    g700(.A(new_n887_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G190gat), .B1(new_n902_), .B2(new_n259_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n611_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n902_), .B2(new_n904_), .ZN(G1351gat));
  NOR2_X1   g704(.A1(new_n554_), .A2(new_n645_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n850_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n604_), .ZN(new_n908_));
  XOR2_X1   g707(.A(new_n908_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n323_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(G204gat), .Z(G1353gat));
  AOI21_X1  g710(.A(new_n292_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT127), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n850_), .A2(new_n906_), .A3(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  XOR2_X1   g714(.A(new_n914_), .B(new_n915_), .Z(G1354gat));
  OAI21_X1  g715(.A(G218gat), .B1(new_n907_), .B2(new_n259_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n255_), .A2(G218gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n907_), .B2(new_n918_), .ZN(G1355gat));
endmodule


