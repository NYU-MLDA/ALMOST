//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(KEYINPUT22), .B1(new_n202_), .B2(KEYINPUT77), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT77), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT78), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT23), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n211_), .B(new_n213_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n218_), .B1(G183gat), .B2(G190gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  OR3_X1    g024(.A1(new_n225_), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT26), .B(G190gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT25), .B1(new_n225_), .B2(KEYINPUT75), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n202_), .A2(new_n207_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n230_), .A2(KEYINPUT24), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OR3_X1    g032(.A1(new_n224_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n222_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT30), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n235_), .B(KEYINPUT30), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT80), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT79), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G15gat), .B(G43gat), .Z(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n242_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n239_), .A2(new_n248_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G113gat), .B(G120gat), .Z(new_n252_));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT82), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n254_), .B(new_n256_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n250_), .A2(new_n251_), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G228gat), .ZN(new_n261_));
  INV_X1    g060(.A(G233gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT88), .B(G211gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G218gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(G197gat), .B(G204gat), .Z(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(KEYINPUT89), .A3(KEYINPUT21), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(KEYINPUT21), .B2(new_n266_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(new_n265_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT83), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n273_), .B2(KEYINPUT1), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(KEYINPUT84), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(KEYINPUT84), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT2), .ZN(new_n287_));
  OAI22_X1  g086(.A1(new_n280_), .A2(new_n286_), .B1(new_n278_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(new_n286_), .B2(new_n280_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n279_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n289_), .B1(new_n290_), .B2(KEYINPUT2), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n275_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n285_), .A2(new_n292_), .ZN(new_n293_));
  AOI211_X1 g092(.A(new_n263_), .B(new_n272_), .C1(new_n293_), .C2(KEYINPUT29), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n296_));
  INV_X1    g095(.A(KEYINPUT91), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n271_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G218gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n264_), .B(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n300_), .B(new_n267_), .C1(KEYINPUT21), .C2(new_n266_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT91), .A3(new_n269_), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n293_), .A2(new_n296_), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n263_), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n303_), .A2(KEYINPUT92), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT92), .ZN(new_n306_));
  INV_X1    g105(.A(new_n302_), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT91), .B1(new_n301_), .B2(new_n269_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n283_), .A2(new_n284_), .B1(new_n275_), .B2(new_n291_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n296_), .ZN(new_n310_));
  OAI22_X1  g109(.A1(new_n307_), .A2(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n306_), .B1(new_n311_), .B2(new_n263_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n295_), .B1(new_n305_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G78gat), .B(G106gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT92), .B1(new_n303_), .B2(new_n304_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(new_n306_), .A3(new_n263_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n314_), .B(KEYINPUT93), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(new_n295_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G22gat), .B(G50gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT86), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n309_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n309_), .B2(new_n323_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n322_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(new_n321_), .A3(new_n326_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n315_), .A2(new_n320_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(KEYINPUT87), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT87), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n329_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n319_), .B1(new_n318_), .B2(new_n295_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n319_), .ZN(new_n339_));
  AOI211_X1 g138(.A(new_n339_), .B(new_n294_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n337_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(KEYINPUT94), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT94), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n313_), .A2(new_n339_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n320_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n345_), .B2(new_n337_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n260_), .B(new_n333_), .C1(new_n342_), .C2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n293_), .A2(new_n254_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n254_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n309_), .A2(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n348_), .A2(KEYINPUT4), .A3(new_n350_), .ZN(new_n355_));
  OR3_X1    g154(.A1(new_n309_), .A2(KEYINPUT4), .A3(new_n349_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n352_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT0), .ZN(new_n359_));
  INV_X1    g158(.A(G57gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G85gat), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n354_), .A2(new_n357_), .A3(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n362_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n365_), .B(KEYINPUT95), .Z(new_n366_));
  XOR2_X1   g165(.A(new_n366_), .B(KEYINPUT19), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT25), .B(G183gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT96), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n227_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n217_), .A2(new_n219_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n224_), .A2(new_n221_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G169gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n207_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n210_), .ZN(new_n379_));
  OAI22_X1  g178(.A1(new_n374_), .A2(new_n375_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n369_), .B1(new_n380_), .B2(new_n271_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n272_), .A2(new_n222_), .A3(new_n234_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n368_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n380_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n367_), .B1(new_n385_), .B2(new_n272_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n369_), .B1(new_n235_), .B2(new_n271_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT32), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n384_), .A2(new_n388_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT99), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT99), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n384_), .A2(new_n397_), .A3(new_n388_), .A4(new_n394_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n363_), .A2(new_n364_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT101), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n381_), .A2(new_n382_), .A3(new_n368_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n385_), .A2(new_n298_), .A3(new_n302_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n368_), .B1(new_n402_), .B2(new_n387_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n403_), .B2(KEYINPUT100), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n403_), .A2(KEYINPUT100), .ZN(new_n405_));
  OAI211_X1 g204(.A(KEYINPUT32), .B(new_n393_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n399_), .A2(new_n400_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n400_), .B1(new_n399_), .B2(new_n406_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n393_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n386_), .A2(new_n387_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(new_n383_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n384_), .A2(new_n393_), .A3(new_n388_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n355_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n362_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n364_), .A2(KEYINPUT33), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n419_), .B(new_n362_), .C1(new_n354_), .C2(new_n357_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT98), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n417_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n347_), .B1(new_n409_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n333_), .B1(new_n342_), .B2(new_n346_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n410_), .B1(new_n405_), .B2(new_n404_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n413_), .A2(KEYINPUT27), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT27), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n414_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n427_), .A2(new_n260_), .A3(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n430_), .A2(KEYINPUT102), .A3(new_n432_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT102), .B1(new_n430_), .B2(new_n432_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n333_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n341_), .A2(KEYINPUT94), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n345_), .A2(new_n343_), .A3(new_n337_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n260_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n437_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n434_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n363_), .A2(new_n364_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n426_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G29gat), .B(G36gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G43gat), .B(G50gat), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n449_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT15), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455_));
  INV_X1    g254(.A(G1gat), .ZN(new_n456_));
  INV_X1    g255(.A(G8gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G8gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT15), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n452_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n454_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G229gat), .A2(G233gat), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n453_), .A2(new_n461_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT72), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT72), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n464_), .A2(new_n469_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n461_), .B(new_n453_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(G229gat), .A3(G233gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n468_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G113gat), .B(G141gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G197gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT73), .B(G169gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n468_), .A2(new_n472_), .A3(new_n470_), .A4(new_n477_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT74), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n480_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT74), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n447_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT70), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT71), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  AND2_X1   g292(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT64), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT64), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n493_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT65), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G85gat), .A2(G92gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G85gat), .A2(G92gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT9), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(G85gat), .A3(G92gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n501_), .A2(new_n502_), .A3(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n498_), .A2(KEYINPUT64), .A3(new_n499_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n496_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n517_));
  AOI21_X1  g316(.A(G106gat), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(G85gat), .A2(G92gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(KEYINPUT9), .A3(new_n503_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n523_), .A3(new_n511_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT65), .B1(new_n518_), .B2(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n515_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527_));
  INV_X1    g326(.A(G99gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(new_n493_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n510_), .A2(new_n512_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n504_), .A2(new_n505_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT8), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n530_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT66), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT66), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n529_), .A2(new_n541_), .A3(new_n530_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n521_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n534_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n537_), .B1(new_n544_), .B2(KEYINPUT8), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n463_), .B(new_n454_), .C1(new_n526_), .C2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT34), .ZN(new_n548_));
  INV_X1    g347(.A(new_n534_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n532_), .B1(new_n531_), .B2(KEYINPUT66), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(new_n542_), .ZN(new_n551_));
  OAI22_X1  g350(.A1(new_n551_), .A2(new_n535_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n515_), .A2(new_n525_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI221_X1 g353(.A(new_n546_), .B1(KEYINPUT35), .B2(new_n548_), .C1(new_n453_), .C2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(KEYINPUT35), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(KEYINPUT36), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n556_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n555_), .B(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n560_), .B(KEYINPUT36), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n489_), .A2(KEYINPUT70), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n492_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n562_), .A2(new_n566_), .A3(new_n570_), .A4(new_n491_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(new_n225_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(G211gat), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n461_), .B(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G71gat), .B(G78gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n581_), .B1(KEYINPUT11), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n580_), .B(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n578_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n576_), .A2(new_n577_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n578_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n572_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G120gat), .B(G148gat), .ZN(new_n593_));
  INV_X1    g392(.A(G204gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT5), .B(G176gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G230gat), .A2(G233gat), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n583_), .B(new_n584_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n526_), .A2(new_n545_), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n585_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT67), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(KEYINPUT67), .B(new_n600_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(KEYINPUT68), .A2(KEYINPUT12), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n601_), .B1(new_n526_), .B2(new_n545_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n552_), .A2(new_n585_), .A3(new_n553_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n609_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(KEYINPUT68), .A2(KEYINPUT12), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n609_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n554_), .B2(new_n601_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n612_), .A2(new_n600_), .A3(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n598_), .B1(new_n608_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n609_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n610_), .B1(new_n613_), .B2(new_n609_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(new_n599_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n621_), .A2(new_n606_), .A3(new_n607_), .A4(new_n597_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT69), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n624_), .B2(KEYINPUT13), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n626_));
  NAND3_X1  g425(.A1(new_n617_), .A2(new_n622_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n592_), .A2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n488_), .A2(new_n456_), .A3(new_n445_), .A4(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n628_), .A2(new_n483_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n590_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n445_), .B1(new_n434_), .B2(new_n443_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n567_), .B(new_n635_), .C1(new_n636_), .C2(new_n426_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G1gat), .B1(new_n637_), .B2(new_n446_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n631_), .A2(new_n632_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n633_), .A2(new_n638_), .A3(new_n639_), .ZN(G1324gat));
  OAI21_X1  g439(.A(G8gat), .B1(new_n637_), .B2(new_n437_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT39), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n643_), .B(G8gat), .C1(new_n637_), .C2(new_n437_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n437_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n488_), .A2(new_n457_), .A3(new_n646_), .A4(new_n630_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT103), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n650_), .A3(new_n647_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n649_), .A2(KEYINPUT40), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT40), .B1(new_n649_), .B2(new_n651_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n637_), .B2(new_n260_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT41), .Z(new_n656_));
  NOR2_X1   g455(.A1(new_n260_), .A2(G15gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n488_), .A2(new_n630_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1326gat));
  XNOR2_X1  g458(.A(new_n441_), .B(KEYINPUT104), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(G22gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n488_), .A2(new_n630_), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G22gat), .B1(new_n637_), .B2(new_n660_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT105), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n665_), .B(G22gat), .C1(new_n637_), .C2(new_n660_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n664_), .A2(KEYINPUT42), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT42), .B1(new_n664_), .B2(new_n666_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n662_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT106), .ZN(G1327gat));
  NOR3_X1   g469(.A1(new_n629_), .A2(new_n591_), .A3(new_n567_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n488_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G29gat), .B1(new_n673_), .B2(new_n445_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT43), .B1(new_n447_), .B2(new_n572_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  INV_X1    g475(.A(new_n572_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n676_), .B(new_n677_), .C1(new_n636_), .C2(new_n426_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n634_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n679_), .A2(KEYINPUT44), .A3(new_n590_), .A4(new_n680_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(G29gat), .A3(new_n445_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n679_), .A2(new_n590_), .A3(new_n680_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n674_), .B1(new_n682_), .B2(new_n685_), .ZN(G1328gat));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  INV_X1    g486(.A(G36gat), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n591_), .B(new_n634_), .C1(new_n675_), .C2(new_n678_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n437_), .B1(new_n689_), .B2(KEYINPUT44), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n690_), .B2(new_n685_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n437_), .A2(G36gat), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n693_));
  NAND3_X1  g492(.A1(new_n673_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n693_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n692_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n672_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n694_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n687_), .B1(new_n691_), .B2(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n689_), .A2(KEYINPUT44), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n681_), .A2(new_n646_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G36gat), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n702_), .A2(KEYINPUT46), .A3(new_n694_), .A4(new_n697_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n699_), .A2(new_n703_), .ZN(G1329gat));
  INV_X1    g503(.A(G43gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(new_n672_), .B2(new_n260_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n681_), .A2(G43gat), .A3(new_n442_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(new_n700_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g508(.A(new_n660_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G50gat), .B1(new_n673_), .B2(new_n710_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n681_), .A2(G50gat), .A3(new_n427_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(new_n685_), .ZN(G1331gat));
  INV_X1    g512(.A(new_n447_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n482_), .A2(new_n591_), .A3(new_n485_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n714_), .A2(new_n629_), .A3(new_n567_), .A4(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n446_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n628_), .A2(new_n483_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n592_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n714_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n445_), .A2(new_n360_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n718_), .B1(new_n722_), .B2(new_n723_), .ZN(G1332gat));
  OAI21_X1  g523(.A(G64gat), .B1(new_n717_), .B2(new_n437_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT48), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n437_), .A2(G64gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n722_), .B2(new_n727_), .ZN(G1333gat));
  OAI21_X1  g527(.A(G71gat), .B1(new_n717_), .B2(new_n260_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT49), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n260_), .A2(G71gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n722_), .B2(new_n731_), .ZN(G1334gat));
  OAI21_X1  g531(.A(G78gat), .B1(new_n717_), .B2(new_n660_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT50), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n660_), .A2(G78gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n722_), .B2(new_n735_), .ZN(G1335gat));
  INV_X1    g535(.A(new_n567_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n720_), .A2(new_n591_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n714_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT108), .ZN(new_n740_));
  AOI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n445_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n679_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n675_), .A2(KEYINPUT109), .A3(new_n678_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n738_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n445_), .A2(G85gat), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT110), .Z(new_n747_));
  AOI21_X1  g546(.A(new_n741_), .B1(new_n745_), .B2(new_n747_), .ZN(G1336gat));
  INV_X1    g547(.A(G92gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n740_), .A2(new_n749_), .A3(new_n646_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n745_), .A2(new_n646_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n749_), .ZN(G1337gat));
  OAI211_X1 g551(.A(new_n740_), .B(new_n442_), .C1(new_n497_), .C2(new_n500_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n743_), .A2(new_n442_), .A3(new_n738_), .A4(new_n744_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G99gat), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT51), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n753_), .A2(new_n755_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1338gat));
  NAND3_X1  g559(.A1(new_n740_), .A2(new_n493_), .A3(new_n427_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n679_), .A2(new_n427_), .A3(new_n590_), .A4(new_n719_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G106gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G106gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT53), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n761_), .B(new_n768_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1339gat));
  AOI21_X1  g569(.A(new_n477_), .B1(new_n471_), .B2(new_n465_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n464_), .A2(new_n466_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n465_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n480_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT112), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n480_), .A2(new_n773_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n622_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n599_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n621_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NOR4_X1   g581(.A1(new_n612_), .A2(new_n615_), .A3(new_n781_), .A4(new_n600_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT56), .B1(new_n785_), .B2(new_n598_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n779_), .B1(new_n786_), .B2(KEYINPUT114), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n600_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n616_), .B1(KEYINPUT55), .B2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n598_), .B1(new_n789_), .B2(new_n783_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n598_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n787_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT115), .B1(new_n798_), .B2(KEYINPUT58), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n787_), .B2(new_n795_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n572_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n483_), .A2(new_n622_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n791_), .B(new_n597_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n786_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n623_), .A2(new_n778_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n737_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT57), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n806_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n810_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n567_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(KEYINPUT113), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n813_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n590_), .B1(new_n805_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n715_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT111), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n572_), .B1(new_n821_), .B2(KEYINPUT111), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT54), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n629_), .B2(new_n715_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n572_), .A4(new_n822_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n825_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n820_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n811_), .A2(new_n812_), .A3(KEYINPUT57), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n817_), .B1(new_n816_), .B2(KEYINPUT113), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT58), .B1(new_n797_), .B2(new_n798_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n677_), .B1(new_n837_), .B2(new_n803_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n591_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT117), .B1(new_n839_), .B2(new_n830_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n833_), .A2(new_n840_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n443_), .A2(new_n446_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n842_), .A2(KEYINPUT118), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(KEYINPUT118), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(G113gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n483_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n841_), .B2(new_n845_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n820_), .A2(new_n831_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n852_), .A2(new_n845_), .A3(KEYINPUT119), .A4(new_n850_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n839_), .A2(new_n830_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n843_), .A2(new_n850_), .A3(new_n844_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n851_), .A2(new_n858_), .A3(new_n487_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n849_), .B1(new_n859_), .B2(new_n848_), .ZN(G1340gat));
  INV_X1    g659(.A(G120gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n628_), .B2(KEYINPUT60), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n847_), .B(new_n862_), .C1(KEYINPUT60), .C2(new_n861_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n851_), .A2(new_n858_), .A3(new_n628_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n861_), .ZN(G1341gat));
  INV_X1    g664(.A(G127gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n846_), .B2(new_n590_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(KEYINPUT120), .B(new_n866_), .C1(new_n846_), .C2(new_n590_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n851_), .A2(new_n858_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n590_), .A2(new_n866_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n869_), .A2(new_n870_), .B1(new_n871_), .B2(new_n872_), .ZN(G1342gat));
  INV_X1    g672(.A(G134gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n847_), .A2(new_n874_), .A3(new_n737_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n851_), .A2(new_n858_), .A3(new_n572_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n874_), .ZN(G1343gat));
  NAND2_X1  g676(.A1(new_n427_), .A2(new_n260_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n878_), .A2(new_n646_), .A3(new_n446_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT121), .Z(new_n880_));
  AND2_X1   g679(.A1(new_n841_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n483_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT122), .B(G141gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n881_), .A2(new_n629_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n591_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  INV_X1    g688(.A(G162gat), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n841_), .A2(new_n890_), .A3(new_n737_), .A4(new_n880_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n841_), .A2(new_n677_), .A3(new_n880_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n890_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  OAI211_X1 g694(.A(KEYINPUT123), .B(new_n891_), .C1(new_n892_), .C2(new_n890_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n437_), .A2(new_n445_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n442_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n852_), .A2(new_n660_), .A3(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901_), .B2(new_n481_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT124), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n904_), .B(G169gat), .C1(new_n901_), .C2(new_n481_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(KEYINPUT62), .A3(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n901_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(new_n377_), .A3(new_n483_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n906_), .B(new_n908_), .C1(KEYINPUT62), .C2(new_n903_), .ZN(G1348gat));
  OAI21_X1  g708(.A(new_n207_), .B1(new_n901_), .B2(new_n628_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n911_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n427_), .B1(new_n833_), .B2(new_n840_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n899_), .A2(new_n207_), .A3(new_n628_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n912_), .A2(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  NOR2_X1   g715(.A1(new_n899_), .A2(new_n590_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n852_), .A2(new_n372_), .A3(new_n660_), .A4(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n914_), .A2(new_n917_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n225_), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n901_), .B2(new_n572_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n737_), .A2(new_n227_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n901_), .B2(new_n923_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(KEYINPUT126), .ZN(G1351gat));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n878_), .A2(new_n445_), .A3(new_n437_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n841_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n926_), .B1(new_n841_), .B2(new_n927_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n483_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(G197gat), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n832_), .B1(new_n820_), .B2(new_n831_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n839_), .A2(KEYINPUT117), .A3(new_n830_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n927_), .B1(new_n933_), .B2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT127), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n928_), .ZN(new_n937_));
  INV_X1    g736(.A(G197gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n937_), .A2(new_n938_), .A3(new_n483_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n932_), .A2(new_n939_), .ZN(G1352gat));
  AOI21_X1  g739(.A(G204gat), .B1(new_n937_), .B2(new_n629_), .ZN(new_n941_));
  AOI211_X1 g740(.A(new_n594_), .B(new_n628_), .C1(new_n936_), .C2(new_n928_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1353gat));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n590_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n937_), .B2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n946_), .ZN(new_n948_));
  AOI211_X1 g747(.A(new_n944_), .B(new_n948_), .C1(new_n936_), .C2(new_n928_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n947_), .A2(new_n949_), .ZN(G1354gat));
  NAND3_X1  g749(.A1(new_n937_), .A2(new_n299_), .A3(new_n737_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n572_), .B1(new_n936_), .B2(new_n928_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n299_), .B2(new_n952_), .ZN(G1355gat));
endmodule


