//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT21), .ZN(new_n202_));
  INV_X1    g001(.A(G197gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  AND3_X1   g004(.A1(new_n205_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT87), .B1(new_n205_), .B2(G197gat), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n202_), .B(new_n204_), .C1(new_n206_), .C2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT88), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT87), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(new_n203_), .B2(G204gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n205_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n213_));
  AOI22_X1  g012(.A1(new_n212_), .A2(new_n213_), .B1(new_n203_), .B2(G204gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(KEYINPUT88), .A3(new_n202_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G211gat), .B(G218gat), .Z(new_n216_));
  INV_X1    g015(.A(KEYINPUT86), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(new_n205_), .B2(G197gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n205_), .A2(G197gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n203_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n216_), .B1(new_n221_), .B2(KEYINPUT21), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n210_), .A2(new_n215_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT89), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT89), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n210_), .A2(new_n215_), .A3(new_n222_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n216_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n228_), .A2(new_n214_), .A3(new_n202_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G169gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT22), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT22), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G169gat), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT82), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT81), .B1(G183gat), .B2(G190gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT23), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n243_), .B(new_n246_), .C1(G183gat), .C2(G190gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n236_), .A2(KEYINPUT82), .A3(new_n237_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n240_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G190gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT26), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT26), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G190gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G183gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT25), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G183gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n245_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n244_), .A2(KEYINPUT23), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT80), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n265_), .A2(KEYINPUT24), .A3(new_n237_), .A4(new_n266_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n260_), .A2(new_n263_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n249_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n227_), .A2(new_n230_), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n229_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n257_), .A2(new_n259_), .A3(KEYINPUT90), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT90), .B1(new_n257_), .B2(new_n259_), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n254_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n268_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n270_), .A2(new_n243_), .A3(new_n246_), .A4(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n261_), .A2(new_n262_), .B1(new_n256_), .B2(new_n250_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n237_), .B(KEYINPUT91), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n236_), .ZN(new_n283_));
  OAI22_X1  g082(.A1(new_n278_), .A2(new_n280_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n274_), .B(KEYINPUT20), .C1(new_n275_), .C2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G226gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT19), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n227_), .A2(new_n230_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n289_), .B2(new_n272_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT20), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n275_), .B2(new_n285_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n286_), .A2(new_n288_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G8gat), .B(G36gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT18), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G64gat), .ZN(new_n296_));
  INV_X1    g095(.A(G92gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT20), .B1(new_n275_), .B2(new_n285_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n227_), .A2(new_n230_), .A3(new_n273_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n300_), .A2(new_n301_), .A3(new_n288_), .ZN(new_n302_));
  AOI211_X1 g101(.A(new_n229_), .B(new_n284_), .C1(new_n224_), .C2(new_n226_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT94), .B1(new_n303_), .B2(new_n291_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT94), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n305_), .B(KEYINPUT20), .C1(new_n289_), .C2(new_n284_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n289_), .A2(new_n272_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n302_), .B1(new_n308_), .B2(new_n288_), .ZN(new_n309_));
  OAI211_X1 g108(.A(KEYINPUT27), .B(new_n299_), .C1(new_n309_), .C2(new_n298_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n288_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n290_), .A2(new_n292_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n298_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n298_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n311_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT84), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT1), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n318_), .B(new_n320_), .C1(new_n323_), .C2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n321_), .B(KEYINPUT84), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n319_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n318_), .B(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n327_), .B(new_n324_), .C1(new_n329_), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT85), .B1(new_n333_), .B2(KEYINPUT29), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n289_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G78gat), .B(G106gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G22gat), .B(G50gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(KEYINPUT28), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n333_), .B2(KEYINPUT29), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G228gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n339_), .A2(new_n326_), .A3(new_n332_), .A4(new_n343_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n342_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n336_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n289_), .A2(new_n348_), .A3(new_n334_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n337_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n347_), .B1(new_n337_), .B2(new_n349_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G127gat), .B(G134gat), .Z(new_n354_));
  XOR2_X1   g153(.A(G113gat), .B(G120gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n333_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n326_), .A3(new_n332_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT92), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G1gat), .B(G29gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT0), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G57gat), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n364_), .A2(KEYINPUT0), .ZN(new_n367_));
  INV_X1    g166(.A(G57gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(KEYINPUT0), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n366_), .A2(new_n370_), .A3(G85gat), .ZN(new_n371_));
  AOI21_X1  g170(.A(G85gat), .B1(new_n366_), .B2(new_n370_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n358_), .A2(KEYINPUT4), .A3(new_n359_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n333_), .A2(new_n357_), .A3(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n362_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n363_), .B(new_n373_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n360_), .A2(new_n362_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n381_));
  OAI22_X1  g180(.A1(new_n380_), .A2(new_n381_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n272_), .B(KEYINPUT30), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G15gat), .B(G43gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n272_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n387_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n385_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n388_), .A2(new_n392_), .A3(new_n385_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT31), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT83), .B1(new_n356_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n396_), .B2(new_n356_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(new_n395_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n395_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n403_), .B2(new_n393_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  NOR4_X1   g204(.A1(new_n317_), .A2(new_n353_), .A3(new_n383_), .A4(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n315_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n382_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n358_), .A2(new_n362_), .A3(new_n359_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n373_), .A2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n382_), .B2(new_n408_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n407_), .A2(new_n409_), .A3(new_n299_), .A4(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT93), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n298_), .A2(KEYINPUT32), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n293_), .B2(new_n416_), .ZN(new_n417_));
  AND4_X1   g216(.A1(new_n415_), .A2(new_n312_), .A3(new_n313_), .A4(new_n416_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n383_), .B1(new_n309_), .B2(new_n416_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n414_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n352_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n383_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n310_), .A2(KEYINPUT96), .A3(new_n316_), .A4(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n310_), .A2(new_n316_), .A3(new_n423_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n422_), .A2(new_n424_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n406_), .B1(new_n428_), .B2(new_n405_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G71gat), .B(G78gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G57gat), .B(G64gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT11), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n431_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(KEYINPUT11), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(new_n431_), .A3(KEYINPUT11), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT69), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT7), .ZN(new_n442_));
  INV_X1    g241(.A(G99gat), .ZN(new_n443_));
  INV_X1    g242(.A(G106gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G99gat), .A2(G106gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n445_), .A2(new_n448_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT65), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT8), .ZN(new_n453_));
  XOR2_X1   g252(.A(G85gat), .B(G92gat), .Z(new_n454_));
  NAND3_X1  g253(.A1(new_n451_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n453_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n457_));
  INV_X1    g256(.A(G85gat), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n458_), .A2(KEYINPUT64), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(KEYINPUT64), .ZN(new_n460_));
  OAI21_X1  g259(.A(G92gat), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n458_), .A2(new_n297_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n461_), .A2(new_n462_), .B1(KEYINPUT9), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT10), .B(G99gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n448_), .B(new_n449_), .C1(new_n465_), .C2(G106gat), .ZN(new_n466_));
  OAI22_X1  g265(.A1(new_n456_), .A2(new_n457_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n437_), .A2(KEYINPUT69), .A3(new_n438_), .ZN(new_n468_));
  AND4_X1   g267(.A1(KEYINPUT12), .A2(new_n441_), .A3(new_n467_), .A4(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(KEYINPUT66), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT66), .ZN(new_n471_));
  OAI221_X1 g270(.A(new_n471_), .B1(new_n464_), .B2(new_n466_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n439_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT12), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n469_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n470_), .A2(new_n472_), .A3(new_n439_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT70), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G230gat), .A2(G233gat), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n477_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n439_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n478_), .B1(new_n484_), .B2(KEYINPUT67), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n470_), .A2(new_n472_), .A3(new_n486_), .A4(new_n439_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n480_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT68), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT68), .ZN(new_n491_));
  AOI211_X1 g290(.A(new_n491_), .B(new_n480_), .C1(new_n485_), .C2(new_n487_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n483_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G120gat), .B(G148gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(G204gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT5), .B(G176gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT71), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n483_), .B(new_n497_), .C1(new_n490_), .C2(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT13), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT13), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n503_), .A3(new_n500_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506_));
  INV_X1    g305(.A(G1gat), .ZN(new_n507_));
  INV_X1    g306(.A(G8gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT14), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G1gat), .B(G8gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G29gat), .B(G36gat), .Z(new_n513_));
  XOR2_X1   g312(.A(G43gat), .B(G50gat), .Z(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G29gat), .B(G36gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G43gat), .B(G50gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n512_), .B(new_n519_), .Z(new_n520_));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n515_), .A2(KEYINPUT15), .A3(new_n518_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT15), .B1(new_n515_), .B2(new_n518_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n512_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n512_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n519_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n529_), .A3(new_n521_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(G169gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n203_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n523_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT79), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n534_), .A2(new_n535_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n523_), .A2(new_n530_), .ZN(new_n539_));
  OAI22_X1  g338(.A1(new_n537_), .A2(new_n538_), .B1(new_n539_), .B2(new_n533_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n505_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n470_), .A2(new_n472_), .A3(new_n519_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n526_), .A2(new_n467_), .A3(KEYINPUT73), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT73), .B1(new_n526_), .B2(new_n467_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n543_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT74), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n526_), .A2(new_n467_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n526_), .A2(new_n467_), .A3(KEYINPUT73), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n547_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT35), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n546_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n554_), .A2(KEYINPUT35), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT74), .B1(new_n544_), .B2(new_n545_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n555_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n556_), .B1(new_n560_), .B2(new_n546_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT77), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n556_), .B(KEYINPUT77), .C1(new_n560_), .C2(new_n546_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT36), .Z(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n564_), .A3(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(KEYINPUT36), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n561_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n576_));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G183gat), .B(G211gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n441_), .A2(new_n468_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n512_), .B(new_n584_), .Z(new_n585_));
  AOI21_X1  g384(.A(new_n582_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n585_), .A2(new_n439_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n439_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n580_), .A2(new_n581_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n588_), .A2(new_n582_), .A3(new_n589_), .A4(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n575_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n430_), .A2(new_n542_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n383_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT38), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n505_), .A2(KEYINPUT72), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n502_), .A2(new_n504_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT37), .B1(new_n571_), .B2(new_n573_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n556_), .B(new_n570_), .C1(new_n560_), .C2(new_n546_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n573_), .A2(KEYINPUT37), .A3(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n603_), .A2(new_n592_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n602_), .A2(new_n607_), .A3(new_n541_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n608_), .A2(new_n430_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(new_n507_), .A3(new_n383_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n610_), .A2(KEYINPUT97), .A3(new_n597_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT97), .B1(new_n610_), .B2(new_n597_), .ZN(new_n612_));
  OAI221_X1 g411(.A(new_n596_), .B1(new_n597_), .B2(new_n610_), .C1(new_n611_), .C2(new_n612_), .ZN(G1324gat));
  INV_X1    g412(.A(new_n317_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G8gat), .B1(new_n594_), .B2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(KEYINPUT98), .B(KEYINPUT39), .Z(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n608_), .A2(new_n508_), .A3(new_n317_), .A4(new_n430_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n615_), .A2(KEYINPUT98), .A3(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT99), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n617_), .A2(new_n623_), .A3(new_n618_), .A4(new_n620_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n622_), .A2(KEYINPUT40), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT40), .B1(new_n622_), .B2(new_n624_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1325gat));
  OAI21_X1  g426(.A(G15gat), .B1(new_n594_), .B2(new_n405_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT41), .Z(new_n629_));
  INV_X1    g428(.A(G15gat), .ZN(new_n630_));
  INV_X1    g429(.A(new_n405_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n609_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(G1326gat));
  OAI21_X1  g432(.A(G22gat), .B1(new_n594_), .B2(new_n352_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n609_), .A2(new_n636_), .A3(new_n353_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1327gat));
  NAND2_X1  g437(.A1(new_n542_), .A2(new_n592_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n429_), .A2(new_n574_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n383_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n603_), .A2(new_n605_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT43), .B1(new_n645_), .B2(KEYINPUT100), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n647_), .B1(new_n429_), .B2(new_n645_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n645_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n421_), .A2(new_n352_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n631_), .B1(new_n650_), .B2(new_n424_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n649_), .B(new_n646_), .C1(new_n651_), .C2(new_n406_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n639_), .B1(new_n648_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT44), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(G29gat), .A3(new_n383_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n640_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n644_), .B1(new_n655_), .B2(new_n659_), .ZN(G1328gat));
  NOR3_X1   g459(.A1(new_n642_), .A2(G36gat), .A3(new_n614_), .ZN(new_n661_));
  XOR2_X1   g460(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT103), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n661_), .B(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n614_), .B1(new_n653_), .B2(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n659_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n665_), .B1(new_n667_), .B2(G36gat), .ZN(new_n668_));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT101), .B(new_n669_), .C1(new_n659_), .C2(new_n666_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n664_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT46), .B(new_n664_), .C1(new_n668_), .C2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1329gat));
  INV_X1    g474(.A(KEYINPUT47), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n659_), .A2(G43gat), .A3(new_n631_), .A4(new_n654_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678_));
  INV_X1    g477(.A(G43gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n679_), .B1(new_n642_), .B2(new_n405_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n677_), .A2(new_n678_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n678_), .B1(new_n677_), .B2(new_n680_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n676_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n683_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(KEYINPUT47), .A3(new_n681_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n643_), .B2(new_n353_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n654_), .A2(G50gat), .A3(new_n353_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n659_), .ZN(G1331gat));
  NAND2_X1  g489(.A1(new_n505_), .A2(new_n541_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n429_), .A2(new_n691_), .A3(new_n607_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n368_), .A3(new_n383_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n602_), .A2(new_n541_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n430_), .A2(new_n593_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n694_), .A2(new_n595_), .A3(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n696_), .B2(new_n368_), .ZN(G1332gat));
  INV_X1    g496(.A(G64gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n694_), .A2(new_n695_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n317_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT48), .Z(new_n701_));
  NAND3_X1  g500(.A1(new_n692_), .A2(new_n698_), .A3(new_n317_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1333gat));
  INV_X1    g502(.A(G71gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n699_), .B2(new_n631_), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT105), .B(KEYINPUT49), .Z(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n692_), .A2(new_n704_), .A3(new_n631_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1334gat));
  INV_X1    g508(.A(G78gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n692_), .A2(new_n710_), .A3(new_n353_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n699_), .A2(new_n353_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(G78gat), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n710_), .B(new_n712_), .C1(new_n699_), .C2(new_n353_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(G1335gat));
  INV_X1    g518(.A(new_n592_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n694_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n641_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G85gat), .B1(new_n723_), .B2(new_n383_), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n720_), .B(new_n691_), .C1(new_n648_), .C2(new_n652_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n383_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT108), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n724_), .B1(new_n725_), .B2(new_n727_), .ZN(G1336gat));
  INV_X1    g527(.A(new_n725_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G92gat), .B1(new_n729_), .B2(new_n614_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n317_), .A2(new_n297_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n722_), .B2(new_n731_), .ZN(G1337gat));
  OAI21_X1  g531(.A(G99gat), .B1(new_n729_), .B2(new_n405_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n405_), .A2(new_n465_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n722_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g535(.A1(new_n723_), .A2(new_n444_), .A3(new_n353_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n725_), .A2(new_n353_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G106gat), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT52), .B(new_n444_), .C1(new_n725_), .C2(new_n353_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT109), .B(KEYINPUT53), .Z(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(G1339gat));
  INV_X1    g543(.A(G113gat), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746_));
  INV_X1    g545(.A(new_n538_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n527_), .A2(new_n529_), .A3(new_n522_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n533_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n747_), .A2(new_n536_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n500_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n483_), .A2(new_n752_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n477_), .B(KEYINPUT55), .C1(new_n481_), .C2(new_n482_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n477_), .A2(new_n478_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n489_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(new_n754_), .A3(new_n756_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n498_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT56), .B1(new_n757_), .B2(new_n498_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n746_), .B(new_n751_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT58), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT112), .B1(new_n761_), .B2(KEYINPUT58), .ZN(new_n763_));
  INV_X1    g562(.A(new_n759_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n498_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n763_), .B1(new_n766_), .B2(new_n751_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n649_), .B1(new_n762_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT114), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n500_), .B(new_n540_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n501_), .A2(new_n750_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT57), .B1(new_n772_), .B2(new_n574_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n774_), .B(new_n575_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n649_), .C1(new_n762_), .C2(new_n767_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n592_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n540_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n606_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n599_), .A2(new_n606_), .A3(KEYINPUT110), .A4(new_n541_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT111), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n781_), .A2(KEYINPUT110), .A3(new_n789_), .A4(new_n606_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n786_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT54), .B1(new_n782_), .B2(new_n783_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n790_), .A3(new_n788_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n780_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n317_), .A2(new_n353_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(new_n383_), .A3(new_n631_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n745_), .B1(new_n800_), .B2(new_n541_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n772_), .A2(new_n574_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n774_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n772_), .A2(KEYINPUT57), .A3(new_n574_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n768_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n592_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n794_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n793_), .B1(new_n790_), .B2(new_n788_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n807_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n745_), .A2(KEYINPUT115), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n540_), .A2(G113gat), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(KEYINPUT115), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n798_), .B1(new_n780_), .B2(new_n795_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n812_), .B(new_n815_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n801_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT116), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n801_), .A2(new_n821_), .A3(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1340gat));
  OAI211_X1 g622(.A(new_n812_), .B(new_n602_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT117), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n779_), .A2(new_n592_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT59), .B1(new_n826_), .B2(new_n798_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n602_), .A4(new_n812_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(G120gat), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(G120gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n599_), .B2(KEYINPUT60), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n816_), .B(new_n832_), .C1(KEYINPUT60), .C2(new_n831_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(G1341gat));
  INV_X1    g633(.A(G127gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n800_), .B2(new_n592_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT118), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n835_), .C1(new_n800_), .C2(new_n592_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n827_), .A2(new_n812_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT119), .B(G127gat), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n720_), .A2(new_n842_), .ZN(new_n843_));
  XOR2_X1   g642(.A(new_n843_), .B(KEYINPUT120), .Z(new_n844_));
  AOI22_X1  g643(.A1(new_n837_), .A2(new_n839_), .B1(new_n841_), .B2(new_n844_), .ZN(G1342gat));
  OAI21_X1  g644(.A(G134gat), .B1(new_n840_), .B2(new_n645_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n574_), .A2(G134gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n800_), .B2(new_n847_), .ZN(G1343gat));
  NOR2_X1   g647(.A1(new_n631_), .A2(new_n352_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n850_), .A2(new_n317_), .A3(new_n595_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n796_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n540_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g654(.A(new_n602_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n852_), .A2(new_n856_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT121), .B(G148gat), .Z(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1345gat));
  NOR2_X1   g658(.A1(new_n852_), .A2(new_n592_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT61), .B(G155gat), .Z(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1346gat));
  OR3_X1    g661(.A1(new_n852_), .A2(G162gat), .A3(new_n574_), .ZN(new_n863_));
  OAI21_X1  g662(.A(G162gat), .B1(new_n852_), .B2(new_n645_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1347gat));
  NOR2_X1   g664(.A1(new_n405_), .A2(new_n383_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n317_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n541_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n869_), .A2(KEYINPUT122), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(KEYINPUT122), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n353_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n231_), .B1(new_n810_), .B2(new_n872_), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(KEYINPUT62), .Z(new_n874_));
  AOI211_X1 g673(.A(new_n353_), .B(new_n867_), .C1(new_n795_), .C2(new_n807_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n540_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT123), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n878_), .ZN(G1348gat));
  AOI21_X1  g678(.A(G176gat), .B1(new_n875_), .B2(new_n505_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n826_), .A2(new_n353_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n856_), .A2(new_n235_), .A3(new_n867_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(G1349gat));
  NAND4_X1  g682(.A1(new_n881_), .A2(new_n317_), .A3(new_n866_), .A4(new_n720_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n276_), .A2(new_n277_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n592_), .A2(new_n885_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n884_), .A2(new_n256_), .B1(new_n875_), .B2(new_n886_), .ZN(G1350gat));
  NAND3_X1  g686(.A1(new_n875_), .A2(new_n255_), .A3(new_n575_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n875_), .A2(new_n649_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n250_), .ZN(G1351gat));
  NOR3_X1   g689(.A1(new_n850_), .A2(new_n614_), .A3(new_n383_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n826_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n540_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT124), .B(G197gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1352gat));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n602_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g697(.A(new_n592_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n893_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT125), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n900_), .A2(KEYINPUT126), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(KEYINPUT126), .B1(new_n900_), .B2(new_n902_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n900_), .A2(new_n902_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n903_), .A2(new_n904_), .A3(new_n905_), .ZN(G1354gat));
  INV_X1    g705(.A(G218gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n893_), .A2(new_n907_), .A3(new_n575_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n826_), .A2(new_n645_), .A3(new_n892_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT127), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n908_), .B(new_n912_), .C1(new_n907_), .C2(new_n909_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1355gat));
endmodule


