//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n205_), .B(KEYINPUT88), .Z(new_n206_));
  XOR2_X1   g005(.A(new_n206_), .B(KEYINPUT31), .Z(new_n207_));
  XNOR2_X1  g006(.A(G71gat), .B(G99gat), .ZN(new_n208_));
  INV_X1    g007(.A(G43gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G227gat), .A2(G233gat), .ZN(new_n211_));
  INV_X1    g010(.A(G15gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n210_), .B(new_n213_), .Z(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT86), .B1(new_n217_), .B2(G169gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT22), .B(G169gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n216_), .B(new_n218_), .C1(new_n219_), .C2(KEYINPUT86), .ZN(new_n220_));
  INV_X1    g019(.A(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  OR4_X1    g021(.A1(KEYINPUT87), .A2(new_n221_), .A3(new_n222_), .A4(KEYINPUT23), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT23), .B1(new_n221_), .B2(new_n222_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(KEYINPUT87), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT85), .B(G190gat), .Z(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(G183gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n215_), .B(new_n220_), .C1(new_n228_), .C2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n226_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n215_), .A2(KEYINPUT24), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  MUX2_X1   g033(.A(new_n233_), .B(KEYINPUT24), .S(new_n234_), .Z(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT25), .B(G183gat), .Z(new_n236_));
  NOR2_X1   g035(.A1(new_n222_), .A2(KEYINPUT26), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n229_), .A2(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n232_), .B(new_n235_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n231_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT30), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n231_), .A2(new_n241_), .A3(KEYINPUT30), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n214_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n244_), .A2(new_n214_), .A3(new_n245_), .ZN(new_n247_));
  OR4_X1    g046(.A1(new_n202_), .A2(new_n207_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n248_));
  OR3_X1    g047(.A1(new_n247_), .A2(new_n246_), .A3(new_n202_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n202_), .B1(new_n247_), .B2(new_n246_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n207_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G204gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G197gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n256_), .A2(G197gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT21), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(KEYINPUT95), .B2(new_n257_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(KEYINPUT95), .B2(new_n257_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n260_), .B(new_n261_), .C1(new_n263_), .C2(KEYINPUT21), .ZN(new_n264_));
  INV_X1    g063(.A(new_n261_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(KEYINPUT21), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(KEYINPUT1), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT90), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  OAI211_X1 g071(.A(KEYINPUT90), .B(new_n268_), .C1(new_n269_), .C2(KEYINPUT1), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT91), .B1(new_n268_), .B2(KEYINPUT1), .ZN(new_n274_));
  OR3_X1    g073(.A1(new_n268_), .A2(KEYINPUT91), .A3(KEYINPUT1), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .A4(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G141gat), .ZN(new_n277_));
  INV_X1    g076(.A(G148gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n278_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n276_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n269_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT92), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(KEYINPUT3), .ZN(new_n286_));
  OR3_X1    g085(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n286_), .B(new_n287_), .C1(KEYINPUT2), .C2(new_n279_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n283_), .B(new_n268_), .C1(new_n285_), .C2(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n282_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT29), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n267_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n267_), .A2(KEYINPUT94), .B1(G228gat), .B2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G78gat), .B(G106gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n294_), .A2(new_n296_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n255_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n297_), .A3(new_n254_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n290_), .A2(new_n291_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G22gat), .B(G50gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT96), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n300_), .A2(new_n302_), .A3(new_n307_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n253_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n232_), .B1(G183gat), .B2(G190gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n219_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n312_), .B(new_n215_), .C1(G176gat), .C2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT26), .B(G190gat), .Z(new_n315_));
  OAI21_X1  g114(.A(new_n235_), .B1(new_n236_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n314_), .B1(new_n228_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n267_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n318_), .B(KEYINPUT20), .C1(new_n242_), .C2(new_n267_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT19), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT20), .B1(new_n317_), .B2(new_n267_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n242_), .A2(new_n267_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n321_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT18), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n326_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n330_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT0), .ZN(new_n336_));
  INV_X1    g135(.A(G57gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G85gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n290_), .A2(new_n205_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n206_), .B2(new_n290_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n341_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT98), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  OR3_X1    g148(.A1(new_n206_), .A2(KEYINPUT4), .A3(new_n290_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n342_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT4), .ZN(new_n352_));
  OR3_X1    g151(.A1(new_n345_), .A2(KEYINPUT97), .A3(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT97), .B1(new_n345_), .B2(new_n352_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n331_), .B(new_n334_), .C1(new_n349_), .C2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n346_), .A2(new_n342_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n353_), .A2(new_n354_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n350_), .A2(new_n343_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n341_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT33), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT33), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n364_), .A3(new_n341_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n356_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n361_), .A2(new_n341_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n332_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n319_), .A2(new_n321_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n323_), .A2(KEYINPUT99), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n324_), .B1(new_n323_), .B2(KEYINPUT99), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n321_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n372_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n377_), .A2(new_n369_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n368_), .A2(new_n362_), .B1(new_n370_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n311_), .B1(new_n366_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n310_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n307_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n253_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n252_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n377_), .A2(new_n333_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n386_), .A2(KEYINPUT100), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT100), .B1(new_n386_), .B2(new_n388_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n362_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(new_n367_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n334_), .A2(new_n331_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n387_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n380_), .B1(new_n385_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G230gat), .A2(G233gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n403_));
  INV_X1    g202(.A(G106gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G92gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n339_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G85gat), .A2(G92gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(KEYINPUT9), .A3(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n409_), .A2(KEYINPUT9), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n402_), .A2(new_n406_), .A3(new_n410_), .A4(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT64), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT7), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G99gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n404_), .ZN(new_n418_));
  AND2_X1   g217(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n416_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .A4(new_n404_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n402_), .A3(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n408_), .A2(new_n409_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT8), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT8), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n426_), .A3(new_n423_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n413_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G57gat), .B(G64gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT11), .ZN(new_n430_));
  XOR2_X1   g229(.A(G71gat), .B(G78gat), .Z(new_n431_));
  OR2_X1    g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n429_), .A2(KEYINPUT11), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n431_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n428_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n428_), .A2(new_n435_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n399_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT66), .B(KEYINPUT12), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n412_), .A2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n409_), .A2(KEYINPUT9), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n444_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n445_), .A2(KEYINPUT65), .A3(new_n406_), .A4(new_n410_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n426_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n422_), .A2(new_n426_), .A3(new_n423_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n432_), .B(KEYINPUT12), .C1(new_n433_), .C2(new_n434_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n441_), .A2(new_n398_), .A3(new_n436_), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n439_), .A2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT68), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G120gat), .B(G148gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G176gat), .B(G204gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n457_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n455_), .B(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT13), .Z(new_n463_));
  XNOR2_X1  g262(.A(G113gat), .B(G141gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G169gat), .B(G197gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G43gat), .B(G50gat), .Z(new_n469_));
  INV_X1    g268(.A(G36gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G29gat), .ZN(new_n471_));
  INV_X1    g270(.A(G29gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G36gat), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT69), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT69), .B1(new_n471_), .B2(new_n473_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n469_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT69), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n472_), .A2(G36gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n470_), .A2(G29gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT69), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n476_), .A2(new_n477_), .A3(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G1gat), .B(G8gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT14), .ZN(new_n488_));
  INV_X1    g287(.A(G8gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT78), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT78), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G8gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n488_), .B1(new_n493_), .B2(G1gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n487_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G1gat), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n498_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n495_), .B(new_n486_), .C1(new_n499_), .C2(new_n488_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n477_), .B1(new_n476_), .B2(new_n484_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n485_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n474_), .A2(new_n475_), .A3(new_n469_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n483_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT81), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n476_), .A2(new_n484_), .A3(new_n477_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n506_), .A2(new_n507_), .B1(new_n500_), .B2(new_n497_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n468_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n500_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT78), .B(G8gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n498_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n486_), .B1(new_n512_), .B2(new_n495_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT15), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n476_), .A2(new_n515_), .A3(new_n484_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n476_), .B2(new_n484_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n514_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n501_), .B1(new_n485_), .B2(new_n502_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(KEYINPUT82), .A4(new_n467_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n509_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n467_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT82), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT83), .B1(new_n521_), .B2(new_n524_), .ZN(new_n525_));
  AND4_X1   g324(.A1(KEYINPUT83), .A2(new_n524_), .A3(new_n520_), .A4(new_n509_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n466_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT84), .ZN(new_n528_));
  INV_X1    g327(.A(new_n466_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n521_), .A2(new_n528_), .A3(new_n524_), .A4(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n524_), .A2(new_n520_), .A3(new_n509_), .A4(new_n529_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT84), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n463_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n397_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n450_), .B1(new_n517_), .B2(new_n516_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT35), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT34), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n538_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n476_), .A2(new_n484_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n428_), .A2(KEYINPUT70), .A3(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n412_), .B(new_n544_), .C1(new_n449_), .C2(new_n448_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT70), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n542_), .A2(new_n539_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n543_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n549_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT70), .B1(new_n428_), .B2(new_n544_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n545_), .A2(new_n548_), .A3(KEYINPUT71), .A4(new_n549_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n538_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT72), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n542_), .A2(new_n539_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n559_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n552_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT76), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OAI211_X1 g364(.A(KEYINPUT76), .B(new_n552_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G190gat), .B(G218gat), .Z(new_n567_));
  XOR2_X1   g366(.A(G134gat), .B(G162gat), .Z(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT36), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n565_), .A2(new_n566_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n558_), .A2(new_n560_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT72), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n551_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n576_));
  NAND2_X1  g375(.A1(new_n569_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT74), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n571_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT79), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n435_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n514_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT16), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT17), .B1(new_n585_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT80), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n585_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n590_), .B(new_n592_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n537_), .A2(new_n581_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT103), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n393_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(G1gat), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT75), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n563_), .A2(new_n600_), .A3(new_n570_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n580_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n563_), .B2(new_n570_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT37), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT77), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n571_), .A2(new_n605_), .A3(new_n606_), .A4(new_n580_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n570_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n610_), .A2(new_n566_), .B1(new_n579_), .B2(new_n575_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n605_), .B1(new_n611_), .B2(new_n606_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n593_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n537_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT101), .Z(new_n617_));
  AND3_X1   g416(.A1(new_n617_), .A2(new_n498_), .A3(new_n597_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n617_), .A2(KEYINPUT38), .A3(new_n498_), .A4(new_n597_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(new_n620_), .ZN(new_n622_));
  OAI221_X1 g421(.A(new_n599_), .B1(KEYINPUT38), .B2(new_n618_), .C1(new_n621_), .C2(new_n622_), .ZN(G1324gat));
  NAND2_X1  g422(.A1(new_n391_), .A2(new_n395_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n489_), .B1(new_n594_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT39), .Z(new_n626_));
  NAND3_X1  g425(.A1(new_n617_), .A2(new_n511_), .A3(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(KEYINPUT40), .A3(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1325gat));
  AOI21_X1  g431(.A(new_n212_), .B1(new_n596_), .B2(new_n253_), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n616_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n212_), .A3(new_n253_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1326gat));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n381_), .A2(new_n382_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n596_), .B2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n636_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1327gat));
  NAND2_X1  g444(.A1(new_n397_), .A2(new_n613_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT43), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n397_), .A2(new_n613_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(new_n614_), .A3(new_n536_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n597_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G29gat), .B1(new_n654_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n611_), .A2(new_n614_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n537_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n597_), .A2(new_n472_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT106), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n657_), .B1(new_n661_), .B2(new_n663_), .ZN(G1328gat));
  NAND3_X1  g463(.A1(new_n660_), .A2(new_n470_), .A3(new_n624_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT45), .ZN(new_n666_));
  INV_X1    g465(.A(new_n624_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n653_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n666_), .B1(new_n669_), .B2(new_n470_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT46), .B(new_n666_), .C1(new_n669_), .C2(new_n470_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1329gat));
  OAI21_X1  g473(.A(new_n209_), .B1(new_n661_), .B2(new_n252_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n655_), .A2(G43gat), .A3(new_n253_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n654_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n660_), .B2(new_n640_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n655_), .A2(G50gat), .A3(new_n640_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(new_n653_), .ZN(G1331gat));
  INV_X1    g480(.A(new_n463_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(new_n534_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n615_), .A2(new_n397_), .A3(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n337_), .B1(new_n684_), .B2(new_n393_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n397_), .A2(new_n683_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n686_), .A2(new_n611_), .A3(new_n614_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n597_), .A2(new_n688_), .A3(G57gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n688_), .B2(G57gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n685_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT108), .ZN(G1332gat));
  OR3_X1    g492(.A1(new_n684_), .A2(G64gat), .A3(new_n667_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n687_), .A2(new_n624_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G64gat), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(KEYINPUT48), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(KEYINPUT48), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1333gat));
  NAND2_X1  g498(.A1(new_n687_), .A2(new_n253_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G71gat), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT49), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT49), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n252_), .A2(G71gat), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT109), .ZN(new_n705_));
  OAI22_X1  g504(.A1(new_n702_), .A2(new_n703_), .B1(new_n684_), .B2(new_n705_), .ZN(G1334gat));
  INV_X1    g505(.A(new_n640_), .ZN(new_n707_));
  OR3_X1    g506(.A1(new_n684_), .A2(G78gat), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n687_), .A2(new_n640_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G78gat), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT50), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT50), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(G1335gat));
  NAND2_X1  g512(.A1(new_n683_), .A2(new_n614_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G85gat), .B1(new_n716_), .B2(new_n393_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n686_), .A2(new_n658_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n339_), .A3(new_n597_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1336gat));
  OAI21_X1  g519(.A(G92gat), .B1(new_n716_), .B2(new_n667_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n718_), .A2(new_n407_), .A3(new_n624_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1337gat));
  AOI21_X1  g522(.A(new_n417_), .B1(new_n715_), .B2(new_n253_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n403_), .A2(new_n405_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n253_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT110), .B1(new_n718_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729_));
  NOR4_X1   g528(.A1(new_n686_), .A2(new_n729_), .A3(new_n658_), .A4(new_n726_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n724_), .A2(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT112), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  OAI221_X1 g534(.A(new_n735_), .B1(KEYINPUT111), .B2(KEYINPUT51), .C1(new_n724_), .C2(new_n731_), .ZN(new_n736_));
  AND2_X1   g535(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n734_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1338gat));
  NAND3_X1  g539(.A1(new_n718_), .A2(new_n404_), .A3(new_n640_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n404_), .B1(new_n715_), .B2(new_n640_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n742_), .A2(new_n743_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g546(.A(KEYINPUT121), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT120), .ZN(new_n749_));
  INV_X1    g548(.A(G113gat), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n535_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT59), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n454_), .A2(new_n754_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n450_), .A2(new_n452_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n756_), .A2(KEYINPUT55), .A3(new_n398_), .A4(new_n441_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n453_), .A2(new_n436_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n440_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n412_), .B1(new_n449_), .B2(new_n448_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n435_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n759_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n399_), .B1(new_n758_), .B2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n755_), .A2(new_n757_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n461_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(KEYINPUT56), .A3(new_n461_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n455_), .A2(new_n461_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n527_), .B2(new_n533_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n765_), .A2(KEYINPUT114), .A3(new_n766_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n467_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n518_), .A2(new_n519_), .A3(new_n468_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n466_), .A3(new_n776_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n531_), .A2(KEYINPUT84), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n531_), .A2(KEYINPUT84), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n533_), .A2(KEYINPUT116), .A3(new_n777_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n774_), .A2(KEYINPUT115), .B1(new_n784_), .B2(new_n462_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n770_), .A2(new_n772_), .A3(new_n786_), .A4(new_n773_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n611_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT57), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT77), .B1(new_n581_), .B2(KEYINPUT37), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n771_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n784_), .A2(KEYINPUT58), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT58), .B1(new_n784_), .B2(new_n792_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n791_), .A2(new_n795_), .A3(new_n607_), .A4(new_n604_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n771_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n534_), .A2(new_n797_), .A3(new_n773_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n769_), .A2(new_n768_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n764_), .B2(new_n461_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT115), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n784_), .A2(new_n462_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n787_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n581_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT117), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n790_), .A2(new_n796_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n614_), .ZN(new_n809_));
  OR3_X1    g608(.A1(new_n614_), .A2(KEYINPUT113), .A3(new_n534_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT113), .B1(new_n614_), .B2(new_n534_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n463_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n608_), .B2(new_n612_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT54), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n812_), .C1(new_n608_), .C2(new_n612_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n624_), .B1(new_n809_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n384_), .A2(new_n597_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n753_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n809_), .A2(new_n817_), .ZN(new_n822_));
  XOR2_X1   g621(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n822_), .A2(new_n667_), .A3(new_n820_), .A4(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT119), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n818_), .A2(new_n827_), .A3(new_n820_), .A4(new_n824_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n752_), .B(new_n821_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n818_), .A2(new_n820_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n534_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n748_), .B1(new_n829_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n821_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n752_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n832_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(KEYINPUT121), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n833_), .A2(new_n838_), .ZN(G1340gat));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n840_));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n463_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n831_), .A2(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n834_), .A2(new_n463_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n841_), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n831_), .A2(new_n847_), .A3(new_n593_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n834_), .A2(new_n593_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n831_), .A2(new_n851_), .A3(new_n611_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n834_), .A2(new_n613_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n851_), .ZN(G1343gat));
  NAND2_X1  g653(.A1(new_n383_), .A2(new_n597_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT122), .B1(new_n818_), .B2(new_n856_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n808_), .A2(new_n614_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  NOR4_X1   g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n624_), .A4(new_n855_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n857_), .A2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n535_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n277_), .ZN(G1344gat));
  NOR2_X1   g662(.A1(new_n861_), .A2(new_n682_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(new_n278_), .ZN(G1345gat));
  OAI21_X1  g664(.A(new_n593_), .B1(new_n857_), .B2(new_n860_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT123), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n868_), .B(new_n593_), .C1(new_n857_), .C2(new_n860_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT61), .B(G155gat), .Z(new_n870_));
  AND3_X1   g669(.A1(new_n867_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1346gat));
  INV_X1    g672(.A(new_n613_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G162gat), .B1(new_n861_), .B2(new_n874_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n581_), .A2(G162gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n861_), .B2(new_n876_), .ZN(G1347gat));
  NAND2_X1  g676(.A1(new_n624_), .A2(new_n393_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n878_), .A2(new_n252_), .A3(new_n640_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n822_), .A2(new_n534_), .A3(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n313_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n880_), .A2(G169gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(KEYINPUT62), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(KEYINPUT62), .B2(new_n882_), .ZN(G1348gat));
  NAND2_X1  g683(.A1(new_n822_), .A2(new_n879_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n682_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n216_), .ZN(G1349gat));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n614_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n236_), .B1(new_n889_), .B2(new_n221_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n889_), .A2(G183gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n888_), .B2(new_n892_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n885_), .B2(new_n874_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n581_), .A2(new_n315_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n885_), .B2(new_n895_), .ZN(G1351gat));
  NOR3_X1   g695(.A1(new_n878_), .A2(new_n253_), .A3(new_n707_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n822_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n822_), .A2(KEYINPUT125), .A3(new_n897_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n534_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G197gat), .ZN(G1352gat));
  OAI211_X1 g703(.A(new_n902_), .B(new_n463_), .C1(KEYINPUT126), .C2(new_n256_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n256_), .A2(KEYINPUT126), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1353gat));
  AOI21_X1  g706(.A(new_n614_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  AND2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(new_n908_), .B2(new_n909_), .ZN(G1354gat));
  AOI21_X1  g711(.A(new_n581_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n913_), .A2(KEYINPUT127), .ZN(new_n914_));
  AOI21_X1  g713(.A(G218gat), .B1(new_n913_), .B2(KEYINPUT127), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n613_), .A2(G218gat), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n914_), .A2(new_n915_), .B1(new_n902_), .B2(new_n916_), .ZN(G1355gat));
endmodule


