//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n836_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n202_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT10), .B(G99gat), .Z(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n203_), .A2(new_n204_), .A3(G85gat), .A4(G92gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n207_), .A2(new_n210_), .A3(new_n211_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT7), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n218_), .B(new_n219_), .C1(G99gat), .C2(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n221_), .B(new_n209_), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT70), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n216_), .A2(KEYINPUT69), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT69), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n213_), .A2(new_n215_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT70), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n222_), .A3(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n224_), .A2(new_n225_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n202_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(KEYINPUT71), .A3(KEYINPUT8), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n223_), .A2(new_n216_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT68), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n234_), .A2(KEYINPUT68), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n202_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n234_), .B1(new_n230_), .B2(new_n202_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT71), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n217_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT72), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n217_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n238_), .B1(new_n241_), .B2(KEYINPUT71), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n248_));
  INV_X1    g047(.A(new_n202_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n220_), .A2(new_n222_), .A3(new_n228_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n228_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n227_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n226_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n249_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n248_), .B1(new_n256_), .B2(new_n234_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n246_), .B1(new_n247_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT72), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G57gat), .B(G64gat), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(KEYINPUT11), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(KEYINPUT11), .ZN(new_n262_));
  XOR2_X1   g061(.A(G71gat), .B(G78gat), .Z(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n262_), .A2(new_n263_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT12), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n245_), .A2(new_n259_), .A3(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n266_), .B(new_n217_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G230gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT73), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n258_), .B2(new_n266_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n271_), .A2(new_n279_), .A3(new_n274_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n270_), .A2(new_n276_), .A3(new_n278_), .A4(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n243_), .A2(new_n267_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n271_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n274_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G120gat), .B(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT5), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G176gat), .B(G204gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n290_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n281_), .A2(new_n285_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT13), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT13), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(new_n296_), .A3(new_n293_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(KEYINPUT74), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(KEYINPUT74), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G113gat), .B(G141gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G169gat), .B(G197gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G15gat), .B(G22gat), .ZN(new_n307_));
  INV_X1    g106(.A(G1gat), .ZN(new_n308_));
  INV_X1    g107(.A(G8gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT14), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G1gat), .B(G8gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G29gat), .B(G36gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(G43gat), .B(G50gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G43gat), .B(G50gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(G29gat), .B(G36gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n313_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT15), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n320_), .B(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(new_n323_), .B2(new_n313_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G229gat), .A2(G233gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n313_), .B(new_n320_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n328_), .A2(new_n325_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n306_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT79), .ZN(new_n331_));
  OR3_X1    g130(.A1(new_n327_), .A2(new_n329_), .A3(new_n306_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n302_), .A2(new_n335_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT82), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n337_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  OR3_X1    g142(.A1(new_n343_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT84), .B1(new_n343_), .B2(KEYINPUT23), .ZN(new_n345_));
  INV_X1    g144(.A(new_n343_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n344_), .B(new_n345_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT25), .B(G183gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT26), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT81), .B1(new_n350_), .B2(G190gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G190gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n349_), .B(new_n351_), .C1(new_n352_), .C2(KEYINPUT81), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n342_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT86), .B(G176gat), .ZN(new_n355_));
  INV_X1    g154(.A(G169gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT85), .B1(new_n356_), .B2(KEYINPUT22), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G169gat), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n355_), .B(new_n357_), .C1(new_n358_), .C2(KEYINPUT85), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n343_), .A2(KEYINPUT23), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n359_), .B(new_n339_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n354_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G15gat), .B(G43gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT88), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n369_), .B(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n366_), .B(new_n372_), .Z(new_n373_));
  AND2_X1   g172(.A1(new_n373_), .A2(KEYINPUT89), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(KEYINPUT89), .ZN(new_n375_));
  XOR2_X1   g174(.A(G127gat), .B(G134gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(G113gat), .B(G120gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT31), .Z(new_n379_));
  OR3_X1    g178(.A1(new_n374_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n373_), .A2(KEYINPUT89), .A3(new_n379_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n352_), .A2(new_n349_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n340_), .B1(G169gat), .B2(G176gat), .ZN(new_n385_));
  NOR4_X1   g184(.A1(new_n361_), .A2(new_n384_), .A3(new_n337_), .A4(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n348_), .B1(G183gat), .B2(G190gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n358_), .A2(new_n355_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n388_), .A2(new_n339_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G197gat), .B(G204gat), .Z(new_n391_));
  XNOR2_X1  g190(.A(G211gat), .B(G218gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(KEYINPUT21), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(KEYINPUT21), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT20), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT19), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n395_), .B1(new_n354_), .B2(new_n363_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n397_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(new_n354_), .A3(new_n363_), .ZN(new_n402_));
  OAI211_X1 g201(.A(KEYINPUT20), .B(new_n402_), .C1(new_n390_), .C2(new_n395_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n403_), .A2(new_n399_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G8gat), .B(G36gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT18), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT93), .B1(new_n405_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n405_), .A2(new_n409_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n405_), .A2(KEYINPUT93), .A3(new_n409_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n383_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n403_), .A2(new_n399_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n397_), .A2(KEYINPUT97), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n400_), .B1(new_n397_), .B2(KEYINPUT97), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n416_), .B1(new_n419_), .B2(new_n399_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n409_), .B(KEYINPUT99), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT27), .B(new_n411_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n415_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G155gat), .A2(G162gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(G141gat), .A2(G148gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n427_), .B(KEYINPUT3), .Z(new_n428_));
  NAND2_X1  g227(.A1(G141gat), .A2(G148gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT2), .Z(new_n430_));
  OAI211_X1 g229(.A(new_n424_), .B(new_n426_), .C1(new_n428_), .C2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n425_), .B1(KEYINPUT1), .B2(new_n424_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(KEYINPUT1), .B2(new_n424_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n427_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n429_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n436_), .B(new_n378_), .Z(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT4), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(new_n441_), .A3(new_n378_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n437_), .A2(new_n439_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G29gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G57gat), .B(G85gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n445_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n450_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n436_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT29), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n456_), .A2(KEYINPUT28), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(KEYINPUT28), .ZN(new_n458_));
  XOR2_X1   g257(.A(G22gat), .B(G50gat), .Z(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n460_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT92), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n463_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT92), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n461_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n395_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G228gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n471_), .A2(G228gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(G233gat), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n470_), .A2(new_n476_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G78gat), .B(G106gat), .ZN(new_n479_));
  OR3_X1    g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n479_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT90), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n468_), .A2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n482_), .A2(new_n464_), .A3(new_n467_), .A4(KEYINPUT90), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n423_), .A2(new_n453_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n409_), .A2(KEYINPUT32), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n489_), .B(KEYINPUT96), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n405_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n420_), .A2(new_n489_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT98), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n420_), .A2(KEYINPUT98), .A3(new_n489_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n453_), .B(new_n491_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n414_), .B1(new_n411_), .B2(new_n410_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n445_), .A2(KEYINPUT33), .A3(new_n450_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n450_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT95), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT33), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n452_), .A2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n497_), .A2(new_n498_), .A3(new_n502_), .A4(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n488_), .B1(new_n496_), .B2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n382_), .B1(new_n487_), .B2(new_n506_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n486_), .B(new_n422_), .C1(new_n497_), .C2(KEYINPUT27), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT100), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT100), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n415_), .A2(new_n510_), .A3(new_n486_), .A4(new_n422_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n382_), .A2(new_n453_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n507_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n336_), .A2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G190gat), .B(G218gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(G134gat), .B(G162gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT36), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n245_), .A2(new_n323_), .A3(new_n259_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G232gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT34), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n320_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n258_), .A2(new_n528_), .B1(new_n525_), .B2(new_n524_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n521_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n527_), .B1(new_n521_), .B2(new_n529_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n520_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n530_), .A2(new_n531_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT36), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n519_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT75), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT76), .B1(new_n533_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT76), .ZN(new_n539_));
  NOR4_X1   g338(.A1(new_n530_), .A2(new_n531_), .A3(new_n539_), .A4(new_n536_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n532_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT37), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(KEYINPUT37), .B(new_n532_), .C1(new_n538_), .C2(new_n540_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G127gat), .B(G155gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT16), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT77), .ZN(new_n548_));
  XOR2_X1   g347(.A(G183gat), .B(G211gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT17), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(KEYINPUT17), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n313_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(new_n266_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT78), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT78), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n553_), .A2(new_n556_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n545_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n516_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(new_n308_), .A3(new_n453_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT38), .ZN(new_n566_));
  INV_X1    g365(.A(new_n516_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n541_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(new_n561_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n453_), .ZN(new_n571_));
  OAI21_X1  g370(.A(G1gat), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(G1324gat));
  INV_X1    g372(.A(KEYINPUT101), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n567_), .A2(new_n569_), .A3(new_n423_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(G8gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(new_n576_), .B2(KEYINPUT39), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT39), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n575_), .A2(KEYINPUT101), .A3(new_n578_), .A4(G8gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(KEYINPUT39), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n564_), .A2(new_n309_), .A3(new_n423_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT40), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(G1325gat));
  INV_X1    g384(.A(new_n564_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n586_), .A2(G15gat), .A3(new_n382_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT102), .ZN(new_n588_));
  OAI21_X1  g387(.A(G15gat), .B1(new_n570_), .B2(new_n382_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n589_), .A2(KEYINPUT41), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(KEYINPUT41), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n588_), .A2(new_n590_), .A3(new_n591_), .ZN(G1326gat));
  OAI21_X1  g391(.A(G22gat), .B1(new_n570_), .B2(new_n486_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n594_), .ZN(new_n596_));
  OR3_X1    g395(.A1(new_n586_), .A2(G22gat), .A3(new_n486_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(G1327gat));
  XNOR2_X1  g397(.A(new_n333_), .B(KEYINPUT80), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n301_), .A2(new_n561_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n515_), .A2(new_n545_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT43), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT43), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n515_), .A2(new_n603_), .A3(new_n545_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n600_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT44), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(G29gat), .A3(new_n453_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n605_), .A2(KEYINPUT44), .ZN(new_n608_));
  INV_X1    g407(.A(new_n561_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n541_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n567_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n571_), .ZN(new_n612_));
  OAI22_X1  g411(.A1(new_n607_), .A2(new_n608_), .B1(new_n612_), .B2(G29gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT104), .ZN(G1328gat));
  INV_X1    g413(.A(new_n423_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n611_), .A2(G36gat), .A3(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n608_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n615_), .B1(new_n605_), .B2(KEYINPUT44), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT105), .B1(new_n621_), .B2(G36gat), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT105), .ZN(new_n623_));
  INV_X1    g422(.A(G36gat), .ZN(new_n624_));
  AOI211_X1 g423(.A(new_n623_), .B(new_n624_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n618_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT46), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n618_), .B(KEYINPUT46), .C1(new_n622_), .C2(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1329gat));
  INV_X1    g429(.A(new_n382_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n606_), .A2(G43gat), .A3(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n611_), .A2(new_n382_), .ZN(new_n633_));
  OAI22_X1  g432(.A1(new_n632_), .A2(new_n608_), .B1(new_n633_), .B2(G43gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g434(.A(new_n611_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G50gat), .B1(new_n636_), .B2(new_n488_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n606_), .A2(G50gat), .A3(new_n488_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(new_n619_), .ZN(G1331gat));
  AOI21_X1  g438(.A(new_n599_), .B1(new_n507_), .B2(new_n514_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT107), .Z(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(new_n302_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(KEYINPUT108), .A3(new_n562_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n641_), .A2(new_n302_), .A3(new_n562_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT108), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n571_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G57gat), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n640_), .A2(new_n302_), .A3(new_n569_), .ZN(new_n648_));
  INV_X1    g447(.A(G57gat), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n571_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT109), .ZN(G1332gat));
  OAI21_X1  g451(.A(G64gat), .B1(new_n648_), .B2(new_n615_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT48), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n615_), .A2(G64gat), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT110), .Z(new_n656_));
  OAI21_X1  g455(.A(new_n654_), .B1(new_n644_), .B2(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT111), .Z(G1333gat));
  OAI21_X1  g457(.A(G71gat), .B1(new_n648_), .B2(new_n382_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT49), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n382_), .A2(G71gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n644_), .B2(new_n661_), .ZN(G1334gat));
  OAI21_X1  g461(.A(G78gat), .B1(new_n648_), .B2(new_n486_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT50), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n486_), .A2(G78gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT112), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n644_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT113), .ZN(G1335gat));
  AND2_X1   g467(.A1(new_n642_), .A2(new_n610_), .ZN(new_n669_));
  INV_X1    g468(.A(G85gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n453_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n602_), .A2(new_n604_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n672_), .A2(new_n561_), .A3(new_n335_), .A4(new_n302_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G85gat), .B1(new_n673_), .B2(new_n571_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n674_), .ZN(G1336gat));
  INV_X1    g474(.A(G92gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n669_), .A2(new_n676_), .A3(new_n423_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G92gat), .B1(new_n673_), .B2(new_n615_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1337gat));
  AND2_X1   g478(.A1(new_n631_), .A2(new_n208_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n673_), .A2(new_n382_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n669_), .A2(new_n680_), .B1(new_n681_), .B2(G99gat), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT51), .Z(G1338gat));
  OAI21_X1  g482(.A(G106gat), .B1(new_n673_), .B2(new_n486_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT52), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n669_), .A2(new_n209_), .A3(new_n488_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT53), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT53), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n686_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1339gat));
  INV_X1    g490(.A(KEYINPUT120), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT118), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n631_), .A2(new_n453_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT115), .B1(new_n512_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT115), .ZN(new_n698_));
  AOI211_X1 g497(.A(new_n698_), .B(new_n694_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n293_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n335_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT55), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n281_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT12), .B1(new_n243_), .B2(new_n267_), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n244_), .B(new_n246_), .C1(new_n247_), .C2(new_n257_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n257_), .A2(new_n232_), .A3(new_n239_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT72), .B1(new_n708_), .B2(new_n217_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n706_), .B1(new_n710_), .B2(new_n269_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n271_), .A2(new_n279_), .A3(new_n274_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n279_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n714_), .A3(KEYINPUT55), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT114), .B1(new_n711_), .B2(new_n271_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n270_), .A2(KEYINPUT114), .A3(new_n271_), .A4(new_n278_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n284_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n705_), .B(new_n715_), .C1(new_n716_), .C2(new_n718_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n719_), .A2(KEYINPUT56), .A3(new_n290_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT56), .B1(new_n719_), .B2(new_n290_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n703_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n324_), .A2(new_n326_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n306_), .B1(new_n328_), .B2(new_n325_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n331_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n294_), .A2(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n568_), .B1(new_n722_), .B2(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n726_), .A2(new_n293_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT58), .B(new_n729_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n545_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n716_), .A2(new_n718_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n705_), .A2(new_n715_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n290_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT56), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n719_), .A2(KEYINPUT56), .A3(new_n290_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT58), .B1(new_n738_), .B2(new_n729_), .ZN(new_n739_));
  OAI22_X1  g538(.A1(new_n728_), .A2(KEYINPUT57), .B1(new_n731_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n599_), .A2(new_n293_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n727_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n541_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT57), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n561_), .B1(new_n740_), .B2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n599_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n748_), .A2(new_n543_), .A3(new_n609_), .A4(new_n544_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT54), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n701_), .B1(new_n747_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT59), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT116), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n744_), .A2(new_n745_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n728_), .A2(KEYINPUT57), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n729_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT58), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n545_), .A3(new_n730_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n757_), .A2(new_n758_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n751_), .B1(new_n763_), .B2(new_n561_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n756_), .B(KEYINPUT59), .C1(new_n764_), .C2(new_n701_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n755_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT117), .B1(new_n697_), .B2(new_n700_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n696_), .A2(new_n699_), .A3(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n754_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n770_), .A2(new_n764_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n693_), .B1(new_n766_), .B2(new_n772_), .ZN(new_n773_));
  AOI211_X1 g572(.A(KEYINPUT118), .B(new_n771_), .C1(new_n755_), .C2(new_n765_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n599_), .A2(G113gat), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT119), .Z(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n773_), .A2(new_n774_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n753_), .A2(new_n599_), .ZN(new_n779_));
  INV_X1    g578(.A(G113gat), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n692_), .B1(new_n778_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n766_), .A2(new_n772_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT118), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n766_), .A2(new_n693_), .A3(new_n772_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(new_n776_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT120), .A3(new_n781_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n783_), .A2(new_n788_), .ZN(G1340gat));
  OAI21_X1  g588(.A(G120gat), .B1(new_n784_), .B2(new_n301_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT60), .ZN(new_n791_));
  INV_X1    g590(.A(G120gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n302_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n753_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n790_), .A2(new_n795_), .ZN(G1341gat));
  INV_X1    g595(.A(G127gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n753_), .A2(new_n797_), .A3(new_n609_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n773_), .A2(new_n774_), .A3(new_n561_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n797_), .ZN(G1342gat));
  INV_X1    g599(.A(G134gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n753_), .A2(new_n801_), .A3(new_n568_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n545_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n773_), .A2(new_n774_), .A3(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n804_), .B2(new_n801_), .ZN(G1343gat));
  INV_X1    g604(.A(new_n764_), .ZN(new_n806_));
  NOR4_X1   g605(.A1(new_n423_), .A2(new_n631_), .A3(new_n571_), .A4(new_n486_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n599_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n302_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g612(.A1(new_n808_), .A2(new_n561_), .ZN(new_n814_));
  XOR2_X1   g613(.A(KEYINPUT61), .B(G155gat), .Z(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(G1346gat));
  OAI21_X1  g615(.A(G162gat), .B1(new_n808_), .B2(new_n803_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n541_), .A2(G162gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n808_), .B2(new_n818_), .ZN(G1347gat));
  INV_X1    g618(.A(KEYINPUT62), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n423_), .A2(new_n513_), .A3(new_n486_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n806_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n599_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n820_), .B1(new_n824_), .B2(G169gat), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n825_), .A2(KEYINPUT121), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n820_), .A3(G169gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n825_), .B2(KEYINPUT121), .ZN(new_n828_));
  INV_X1    g627(.A(new_n358_), .ZN(new_n829_));
  OAI22_X1  g628(.A1(new_n826_), .A2(new_n828_), .B1(new_n829_), .B2(new_n824_), .ZN(G1348gat));
  NAND3_X1  g629(.A1(new_n823_), .A2(G176gat), .A3(new_n302_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT123), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n355_), .B1(new_n822_), .B2(new_n301_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT122), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1349gat));
  NOR2_X1   g634(.A1(new_n822_), .A2(new_n561_), .ZN(new_n836_));
  MUX2_X1   g635(.A(G183gat), .B(new_n349_), .S(new_n836_), .Z(G1350gat));
  OAI21_X1  g636(.A(G190gat), .B1(new_n822_), .B2(new_n803_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n568_), .A2(new_n352_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n822_), .B2(new_n839_), .ZN(G1351gat));
  NAND3_X1  g639(.A1(new_n488_), .A2(new_n571_), .A3(new_n382_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n423_), .B1(new_n841_), .B2(KEYINPUT124), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(KEYINPUT124), .B2(new_n841_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n806_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n599_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n302_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G204gat), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT125), .Z(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT126), .B1(new_n847_), .B2(G204gat), .ZN(new_n850_));
  OR3_X1    g649(.A1(new_n847_), .A2(KEYINPUT126), .A3(G204gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(G1353gat));
  INV_X1    g651(.A(new_n844_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n561_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n855_));
  AND2_X1   g654(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n854_), .B2(new_n855_), .ZN(G1354gat));
  OR3_X1    g657(.A1(new_n853_), .A2(G218gat), .A3(new_n541_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G218gat), .B1(new_n853_), .B2(new_n803_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1355gat));
endmodule


