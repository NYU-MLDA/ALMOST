//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n940_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_, new_n954_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT0), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(G57gat), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT83), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT84), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT82), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n212_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT1), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n210_), .A2(KEYINPUT84), .A3(new_n211_), .A4(new_n212_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n215_), .A2(new_n218_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G127gat), .B(G134gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n229_), .A2(new_n230_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n210_), .A2(new_n212_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT86), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT86), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT85), .B1(new_n238_), .B2(new_n235_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n235_), .A2(new_n237_), .B1(new_n239_), .B2(new_n226_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n224_), .B(KEYINPUT2), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n218_), .B(new_n234_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n228_), .A2(new_n233_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n237_), .A2(new_n235_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n239_), .A2(new_n226_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n247_), .A2(new_n241_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n248_), .A2(new_n218_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT80), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(new_n250_), .B2(new_n232_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n244_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT4), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n228_), .A2(new_n243_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n232_), .A2(new_n250_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n233_), .B2(new_n250_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT4), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n207_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n207_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n253_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n206_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n255_), .A2(new_n257_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n264_), .B1(new_n265_), .B2(new_n244_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n261_), .B1(new_n266_), .B2(new_n258_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n262_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n205_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT31), .B(G99gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G15gat), .B(G71gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT75), .ZN(new_n273_));
  INV_X1    g072(.A(G169gat), .ZN(new_n274_));
  INV_X1    g073(.A(G176gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(KEYINPUT24), .A3(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n276_), .A2(new_n277_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT24), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT76), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT76), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(G169gat), .A3(G176gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n280_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n278_), .B1(new_n279_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT23), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT23), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(G183gat), .A3(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G190gat), .ZN(new_n292_));
  OR3_X1    g091(.A1(new_n292_), .A2(KEYINPUT74), .A3(KEYINPUT26), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT25), .B(G183gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT26), .B1(new_n292_), .B2(KEYINPUT74), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n286_), .A2(new_n291_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n282_), .A2(new_n284_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n288_), .A2(new_n290_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT22), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(G169gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT22), .B(G169gat), .ZN(new_n305_));
  OAI211_X1 g104(.A(KEYINPUT78), .B(new_n304_), .C1(new_n305_), .C2(new_n302_), .ZN(new_n306_));
  OR4_X1    g105(.A1(new_n302_), .A2(new_n274_), .A3(KEYINPUT78), .A4(KEYINPUT22), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n301_), .B1(new_n308_), .B2(new_n275_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n272_), .B1(new_n297_), .B2(new_n309_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n298_), .A2(KEYINPUT24), .B1(new_n277_), .B2(new_n276_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n278_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n291_), .B(new_n296_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n272_), .ZN(new_n314_));
  AOI21_X1  g113(.A(G176gat), .B1(new_n306_), .B2(new_n307_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n313_), .B(new_n314_), .C1(new_n315_), .C2(new_n301_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G227gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT30), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT81), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n310_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n319_), .B1(new_n310_), .B2(new_n316_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n271_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n310_), .A2(new_n316_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n319_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n271_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n320_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT79), .B(G43gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n257_), .B(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n323_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n328_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n327_), .B1(new_n326_), .B2(new_n320_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n228_), .A2(new_n337_), .A3(new_n243_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G78gat), .B(G106gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n339_), .B(KEYINPUT89), .Z(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n340_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n228_), .A2(new_n343_), .A3(new_n337_), .A4(new_n243_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n342_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n336_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G204gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(G197gat), .ZN(new_n349_));
  INV_X1    g148(.A(G197gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(G204gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G211gat), .B(G218gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n349_), .A2(new_n351_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT21), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(KEYINPUT88), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n352_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n354_), .B(new_n353_), .C1(new_n360_), .C2(KEYINPUT88), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n255_), .B2(KEYINPUT29), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n363_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n342_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n343_), .B1(new_n249_), .B2(new_n337_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n344_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n367_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n336_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n347_), .A2(new_n366_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n366_), .B1(new_n347_), .B2(new_n373_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n331_), .B(new_n335_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n366_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n345_), .A2(new_n346_), .A3(new_n336_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n372_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n347_), .A2(new_n373_), .A3(new_n366_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n323_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n330_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n380_), .B(new_n381_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n270_), .B1(new_n376_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT18), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G64gat), .ZN(new_n388_));
  INV_X1    g187(.A(G92gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT19), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n359_), .A2(new_n361_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n297_), .B2(new_n309_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n397_));
  INV_X1    g196(.A(new_n300_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n291_), .A2(new_n398_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n305_), .A2(new_n275_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT26), .B(G190gat), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n294_), .A2(new_n401_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n402_));
  AND2_X1   g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n274_), .A2(new_n275_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(new_n280_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n278_), .A2(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n399_), .A2(new_n400_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n397_), .B1(new_n407_), .B2(new_n362_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n394_), .B1(new_n396_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n402_), .A2(new_n406_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n400_), .B(new_n298_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n397_), .B1(new_n395_), .B2(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n313_), .B(new_n362_), .C1(new_n315_), .C2(new_n301_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n394_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n391_), .B(KEYINPUT92), .C1(new_n409_), .C2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n396_), .A2(new_n394_), .A3(new_n408_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT91), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n396_), .A2(KEYINPUT91), .A3(new_n408_), .A4(new_n394_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n413_), .A2(new_n414_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(new_n393_), .ZN(new_n424_));
  AOI211_X1 g223(.A(KEYINPUT90), .B(new_n394_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n420_), .B(new_n421_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n417_), .B1(new_n426_), .B2(new_n391_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n409_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n390_), .B1(new_n428_), .B2(new_n415_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT27), .B1(new_n429_), .B2(KEYINPUT92), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(KEYINPUT93), .B(KEYINPUT27), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n420_), .A2(new_n421_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n423_), .A2(new_n393_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT90), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n423_), .A2(new_n422_), .A3(new_n393_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n438_), .A3(new_n390_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n424_), .A2(new_n425_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n420_), .A2(new_n421_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n391_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n433_), .B1(new_n439_), .B2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n431_), .A2(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(KEYINPUT32), .B(new_n390_), .C1(new_n416_), .C2(new_n409_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n434_), .A2(new_n438_), .A3(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n270_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n269_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n267_), .A2(KEYINPUT33), .A3(new_n205_), .A4(new_n268_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n450_), .A2(new_n439_), .A3(new_n442_), .A4(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n253_), .A2(new_n207_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n254_), .A2(new_n259_), .ZN(new_n454_));
  AOI211_X1 g253(.A(new_n205_), .B(new_n453_), .C1(new_n454_), .C2(new_n207_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n448_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n374_), .A2(new_n375_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n382_), .A2(new_n383_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n385_), .A2(new_n444_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G190gat), .B(G218gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G134gat), .ZN(new_n462_));
  INV_X1    g261(.A(G162gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT36), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n464_), .A2(new_n465_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT15), .ZN(new_n469_));
  INV_X1    g268(.A(G29gat), .ZN(new_n470_));
  INV_X1    g269(.A(G36gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(G43gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G29gat), .A2(G36gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G50gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n473_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n472_), .A2(new_n474_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G43gat), .ZN(new_n481_));
  AOI21_X1  g280(.A(G50gat), .B1(new_n481_), .B2(new_n475_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n469_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n477_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(G50gat), .A3(new_n475_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(KEYINPUT15), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT66), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT9), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G92gat), .ZN(new_n490_));
  AND2_X1   g289(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n389_), .A2(G85gat), .ZN(new_n494_));
  INV_X1    g293(.A(G85gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G92gat), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n489_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n488_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n499_), .A2(new_n489_), .A3(G92gat), .A4(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G85gat), .B(G92gat), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n501_), .B(KEYINPUT66), .C1(new_n489_), .C2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT10), .B(G99gat), .Z(new_n504_));
  INV_X1    g303(.A(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT64), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT64), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT6), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT6), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(G99gat), .A3(G106gat), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n504_), .A2(new_n509_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n498_), .A2(new_n503_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n513_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n517_));
  OR3_X1    g316(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT8), .ZN(new_n520_));
  INV_X1    g319(.A(new_n502_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n515_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n468_), .B1(new_n487_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G232gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT34), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n519_), .A2(new_n521_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT8), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n479_), .A2(new_n482_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n515_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n525_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n528_), .A2(new_n529_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n537_), .A2(new_n538_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n466_), .B(new_n467_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT72), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n539_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n546_), .A2(KEYINPUT72), .A3(new_n466_), .A4(new_n467_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n466_), .B(KEYINPUT70), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n539_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n544_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT37), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(new_n551_), .A3(new_n549_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT73), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT73), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n542_), .A2(new_n549_), .A3(new_n554_), .A4(new_n551_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(KEYINPUT37), .A2(new_n550_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G127gat), .B(G155gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT16), .ZN(new_n558_));
  INV_X1    g357(.A(G183gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G211gat), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G15gat), .B(G22gat), .ZN(new_n564_));
  INV_X1    g363(.A(G1gat), .ZN(new_n565_));
  INV_X1    g364(.A(G8gat), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT14), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G1gat), .B(G8gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT11), .ZN(new_n573_));
  AND2_X1   g372(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n574_));
  NOR2_X1   g373(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n574_), .A2(new_n575_), .A3(G78gat), .ZN(new_n576_));
  INV_X1    g375(.A(G78gat), .ZN(new_n577_));
  OR2_X1    g376(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n573_), .B1(new_n576_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G78gat), .B1(new_n574_), .B2(new_n575_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n583_), .A3(KEYINPUT11), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n584_), .A2(new_n585_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n572_), .B(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n563_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n561_), .B(new_n562_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(new_n589_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n460_), .A2(new_n556_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n570_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n535_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n596_), .A2(new_n535_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n595_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n487_), .A2(new_n570_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n594_), .A3(new_n597_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(new_n274_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n350_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n606_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n588_), .A2(new_n524_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n586_), .A2(new_n587_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n534_), .A3(new_n515_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n612_), .A3(KEYINPUT68), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT68), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n588_), .A2(new_n524_), .A3(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n613_), .A2(new_n615_), .A3(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n610_), .A2(new_n612_), .A3(KEYINPUT12), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n588_), .A2(new_n524_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n615_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n618_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT5), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(G176gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(new_n348_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n627_), .B1(new_n618_), .B2(new_n622_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(KEYINPUT13), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT13), .B1(new_n629_), .B2(new_n630_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT69), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT69), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n593_), .A2(new_n609_), .A3(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n270_), .B(KEYINPUT94), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n565_), .A3(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n542_), .A2(new_n549_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n460_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT96), .ZN(new_n646_));
  INV_X1    g445(.A(new_n592_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n631_), .A2(new_n632_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n609_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n646_), .A2(new_n647_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n270_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n643_), .A2(new_n653_), .ZN(G1324gat));
  INV_X1    g453(.A(new_n444_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n639_), .A2(new_n566_), .A3(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n646_), .A2(new_n647_), .A3(new_n650_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n566_), .B1(new_n657_), .B2(new_n655_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n658_), .A2(new_n659_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n656_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT40), .B(new_n656_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1325gat));
  INV_X1    g466(.A(G15gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n639_), .A2(new_n668_), .A3(new_n458_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n458_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G15gat), .B1(new_n651_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n673_), .A2(KEYINPUT41), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(KEYINPUT41), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n669_), .B1(new_n674_), .B2(new_n675_), .ZN(G1326gat));
  INV_X1    g475(.A(G22gat), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n457_), .B(KEYINPUT98), .Z(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n639_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G22gat), .B1(new_n651_), .B2(new_n678_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT42), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(KEYINPUT42), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n684_), .B2(new_n685_), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n550_), .A2(KEYINPUT37), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n553_), .A2(new_n555_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n460_), .A2(new_n689_), .A3(KEYINPUT43), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n376_), .A2(new_n384_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n444_), .A3(new_n652_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n456_), .A2(new_n459_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n691_), .B1(new_n695_), .B2(new_n556_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n592_), .B(new_n650_), .C1(new_n690_), .C2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n698_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(G29gat), .A3(new_n640_), .A4(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n644_), .A2(new_n592_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n695_), .A2(new_n650_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n470_), .B1(new_n705_), .B2(new_n652_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n701_), .A2(new_n706_), .ZN(G1328gat));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n471_), .A3(new_n655_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT100), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT45), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n699_), .A2(new_n655_), .A3(new_n700_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G36gat), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT101), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n713_), .A2(new_n714_), .A3(new_n717_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n710_), .A2(new_n715_), .A3(new_n716_), .A4(new_n712_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1329gat));
  OAI21_X1  g519(.A(new_n473_), .B1(new_n705_), .B2(new_n670_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n670_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n699_), .A2(G43gat), .A3(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(KEYINPUT102), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(KEYINPUT102), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g526(.A1(new_n699_), .A2(G50gat), .A3(new_n457_), .A4(new_n700_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n477_), .B1(new_n705_), .B2(new_n678_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1331gat));
  AND3_X1   g529(.A1(new_n593_), .A2(new_n649_), .A3(new_n648_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G57gat), .B1(new_n731_), .B2(new_n640_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n592_), .A2(new_n609_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n646_), .A2(new_n637_), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT103), .B(G57gat), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n652_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n732_), .B1(new_n735_), .B2(new_n737_), .ZN(G1332gat));
  INV_X1    g537(.A(G64gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n731_), .A2(new_n739_), .A3(new_n655_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n735_), .B2(new_n655_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n742_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(KEYINPUT48), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT48), .B1(new_n743_), .B2(new_n744_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n740_), .B1(new_n745_), .B2(new_n746_), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n734_), .B2(new_n670_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT49), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n670_), .A2(G71gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT105), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n731_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n734_), .B2(new_n678_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n731_), .A2(new_n577_), .A3(new_n679_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1335gat));
  NOR2_X1   g556(.A1(new_n460_), .A2(new_n609_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n702_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n640_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n495_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT106), .Z(new_n763_));
  NOR3_X1   g562(.A1(new_n633_), .A2(new_n647_), .A3(new_n609_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT43), .B1(new_n460_), .B2(new_n689_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n695_), .A2(new_n691_), .A3(new_n556_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n652_), .A2(new_n492_), .A3(new_n491_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n763_), .B1(new_n768_), .B2(new_n769_), .ZN(G1336gat));
  NOR3_X1   g569(.A1(new_n760_), .A2(G92gat), .A3(new_n444_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n768_), .A2(new_n655_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(G92gat), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT107), .ZN(G1337gat));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n758_), .A2(new_n504_), .A3(new_n458_), .A4(new_n759_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT109), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n778_));
  INV_X1    g577(.A(G99gat), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n778_), .B(new_n779_), .C1(new_n768_), .C2(new_n458_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n458_), .B(new_n764_), .C1(new_n690_), .C2(new_n696_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT108), .B1(new_n781_), .B2(G99gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n777_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(KEYINPUT51), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n783_), .B2(KEYINPUT51), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n788_), .B(new_n777_), .C1(new_n780_), .C2(new_n782_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n670_), .B(new_n765_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n778_), .B1(new_n792_), .B2(new_n779_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n781_), .A2(KEYINPUT108), .A3(G99gat), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n795_), .A2(KEYINPUT111), .A3(new_n788_), .A4(new_n777_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n791_), .A2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n775_), .B1(new_n787_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n791_), .A2(new_n796_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(KEYINPUT112), .C1(new_n786_), .C2(new_n785_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1338gat));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802_));
  INV_X1    g601(.A(new_n768_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n457_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n768_), .A2(KEYINPUT113), .A3(new_n457_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(G106gat), .A3(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT52), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n758_), .A2(new_n509_), .A3(new_n457_), .A4(new_n759_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT53), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(new_n812_), .A3(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1339gat));
  NAND3_X1  g613(.A1(new_n689_), .A2(new_n633_), .A3(new_n733_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT54), .Z(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n619_), .A2(new_n621_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n615_), .A2(KEYINPUT115), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n619_), .A2(new_n621_), .B1(new_n821_), .B2(new_n614_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n822_), .B2(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n818_), .A2(new_n614_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n821_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n622_), .B2(KEYINPUT55), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(KEYINPUT56), .A3(new_n627_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT56), .B1(new_n828_), .B2(new_n627_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n828_), .A2(new_n832_), .A3(KEYINPUT56), .A4(new_n627_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n594_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n601_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n606_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n629_), .A2(new_n607_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n817_), .B1(new_n833_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n556_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n828_), .A2(new_n627_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(KEYINPUT116), .A3(new_n829_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n834_), .A2(new_n838_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT58), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT117), .B1(new_n848_), .B2(new_n689_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n846_), .A2(new_n847_), .A3(KEYINPUT58), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n842_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT118), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n609_), .B(new_n629_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n629_), .A2(new_n630_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n607_), .A3(new_n837_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n644_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT57), .Z(new_n857_));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n842_), .A2(new_n849_), .A3(new_n858_), .A4(new_n850_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n852_), .A2(new_n857_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n816_), .B1(new_n860_), .B2(new_n592_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n761_), .A2(new_n655_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(new_n458_), .A3(new_n804_), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT119), .Z(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT59), .B1(new_n861_), .B2(new_n865_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n867_));
  AOI21_X1  g666(.A(new_n647_), .B1(new_n857_), .B2(new_n851_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n864_), .B(new_n867_), .C1(new_n868_), .C2(new_n816_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n870_));
  INV_X1    g669(.A(G113gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n649_), .B2(new_n871_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n866_), .A2(new_n869_), .A3(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n861_), .A2(new_n865_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G113gat), .B1(new_n874_), .B2(new_n609_), .ZN(new_n875_));
  OAI22_X1  g674(.A1(new_n873_), .A2(new_n875_), .B1(new_n870_), .B2(new_n871_), .ZN(G1340gat));
  NAND3_X1  g675(.A1(new_n866_), .A2(new_n637_), .A3(new_n869_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G120gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n860_), .A2(new_n592_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n816_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n882_), .A2(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n633_), .B2(G120gat), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n881_), .A2(new_n864_), .A3(new_n883_), .A4(new_n884_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n885_), .A2(KEYINPUT122), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(KEYINPUT122), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n878_), .B1(new_n886_), .B2(new_n887_), .ZN(G1341gat));
  AOI21_X1  g687(.A(G127gat), .B1(new_n874_), .B2(new_n647_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n866_), .A2(new_n869_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n647_), .A2(G127gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT123), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n889_), .B1(new_n890_), .B2(new_n892_), .ZN(G1342gat));
  AOI21_X1  g692(.A(G134gat), .B1(new_n874_), .B2(new_n644_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n556_), .A2(G134gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n890_), .B2(new_n895_), .ZN(G1343gat));
  AOI21_X1  g695(.A(new_n384_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(new_n609_), .A3(new_n862_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT124), .B(G141gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1344gat));
  NAND3_X1  g699(.A1(new_n897_), .A2(new_n637_), .A3(new_n862_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g701(.A1(new_n897_), .A2(new_n647_), .A3(new_n862_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  AND2_X1   g704(.A1(new_n897_), .A2(new_n862_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n689_), .A2(new_n463_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n897_), .A2(new_n644_), .A3(new_n862_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n906_), .A2(new_n907_), .B1(new_n908_), .B2(new_n463_), .ZN(G1347gat));
  NOR3_X1   g708(.A1(new_n640_), .A2(new_n444_), .A3(new_n670_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n678_), .B(new_n910_), .C1(new_n868_), .C2(new_n816_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G169gat), .B1(new_n911_), .B2(new_n649_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n911_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n915_), .A2(new_n305_), .A3(new_n609_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n912_), .A2(new_n913_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n916_), .A3(new_n917_), .ZN(G1348gat));
  AOI21_X1  g717(.A(G176gat), .B1(new_n915_), .B2(new_n648_), .ZN(new_n919_));
  NOR4_X1   g718(.A1(new_n861_), .A2(new_n275_), .A3(new_n457_), .A4(new_n638_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n910_), .B2(new_n920_), .ZN(G1349gat));
  NAND2_X1  g720(.A1(new_n910_), .A2(new_n647_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n294_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n678_), .B(new_n923_), .C1(new_n868_), .C2(new_n816_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n457_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n922_), .ZN(new_n927_));
  AOI21_X1  g726(.A(KEYINPUT125), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929_));
  NOR4_X1   g728(.A1(new_n861_), .A2(new_n929_), .A3(new_n457_), .A4(new_n922_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n925_), .B1(new_n931_), .B2(new_n559_), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n915_), .A2(new_n644_), .A3(new_n401_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n915_), .A2(new_n556_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(G190gat), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n934_), .B(G190gat), .C1(new_n911_), .C2(new_n689_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n933_), .B1(new_n936_), .B2(new_n938_), .ZN(G1351gat));
  NAND4_X1  g738(.A1(new_n897_), .A2(new_n652_), .A3(new_n655_), .A4(new_n609_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g740(.A1(new_n897_), .A2(new_n652_), .A3(new_n655_), .A4(new_n637_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g742(.A1(new_n897_), .A2(new_n652_), .A3(new_n647_), .A4(new_n655_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n861_), .A2(new_n270_), .A3(new_n384_), .ZN(new_n947_));
  XOR2_X1   g746(.A(KEYINPUT63), .B(G211gat), .Z(new_n948_));
  NAND4_X1  g747(.A1(new_n947_), .A2(new_n647_), .A3(new_n655_), .A4(new_n948_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n946_), .A2(new_n949_), .ZN(G1354gat));
  AND2_X1   g749(.A1(new_n947_), .A2(new_n655_), .ZN(new_n951_));
  INV_X1    g750(.A(G218gat), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n689_), .A2(new_n952_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n947_), .A2(new_n644_), .A3(new_n655_), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n951_), .A2(new_n953_), .B1(new_n954_), .B2(new_n952_), .ZN(G1355gat));
endmodule


