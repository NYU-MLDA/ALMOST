//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n924_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n955_, new_n957_, new_n959_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G230gat), .A2(G233gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G85gat), .B(G92gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  OR3_X1    g010(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n208_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT8), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n217_), .B(new_n208_), .C1(new_n211_), .C2(new_n214_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n208_), .A2(KEYINPUT9), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT64), .B(G92gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT9), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(G85gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n209_), .B(KEYINPUT6), .ZN(new_n224_));
  OR2_X1    g023(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n220_), .A2(new_n223_), .A3(new_n224_), .A4(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n219_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G64gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G57gat), .ZN(new_n232_));
  INV_X1    g031(.A(G57gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G64gat), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n232_), .A2(new_n234_), .A3(KEYINPUT65), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT65), .B1(new_n232_), .B2(new_n234_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT11), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT66), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n239_), .B(KEYINPUT11), .C1(new_n235_), .C2(new_n236_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n232_), .A2(new_n234_), .A3(KEYINPUT65), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n233_), .A2(G64gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n231_), .A2(G57gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT11), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G71gat), .B(G78gat), .Z(new_n248_));
  NAND4_X1  g047(.A1(new_n238_), .A2(new_n240_), .A3(new_n247_), .A4(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n238_), .A2(new_n240_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n230_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n229_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n238_), .A2(new_n240_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n247_), .A2(new_n248_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n254_), .A2(new_n257_), .A3(new_n249_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n252_), .A2(KEYINPUT12), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n249_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n230_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n207_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n206_), .B1(new_n252_), .B2(new_n258_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n205_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n263_), .A2(new_n264_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n205_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NOR4_X1   g070(.A1(new_n263_), .A2(KEYINPUT67), .A3(new_n264_), .A4(new_n205_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n265_), .B(new_n267_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n265_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n259_), .A2(new_n262_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n206_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n264_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n270_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT67), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n269_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n274_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(KEYINPUT13), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n273_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n285_), .A2(new_n286_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n292_));
  NAND2_X1  g091(.A1(G232gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT35), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G43gat), .B(G50gat), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(KEYINPUT72), .B(new_n296_), .C1(new_n230_), .C2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n301_), .B(KEYINPUT15), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n230_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n294_), .A2(new_n295_), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G190gat), .B(G218gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G134gat), .B(G162gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n312_), .A2(KEYINPUT36), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(KEYINPUT71), .Z(new_n314_));
  NAND3_X1  g113(.A1(new_n308_), .A2(new_n309_), .A3(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n312_), .B(KEYINPUT36), .Z(new_n316_));
  INV_X1    g115(.A(new_n309_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(new_n307_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n320_));
  OR3_X1    g119(.A1(new_n319_), .A2(new_n320_), .A3(KEYINPUT37), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n319_), .B2(KEYINPUT37), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n315_), .A2(KEYINPUT73), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n308_), .A2(new_n324_), .A3(new_n309_), .A4(new_n314_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n325_), .A3(new_n318_), .ZN(new_n326_));
  AOI22_X1  g125(.A1(new_n321_), .A2(new_n322_), .B1(KEYINPUT37), .B2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G1gat), .B(G8gat), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n328_), .A2(KEYINPUT75), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(KEYINPUT75), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G15gat), .B(G22gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G1gat), .A2(G8gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT14), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n335_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G231gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(new_n260_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT17), .ZN(new_n342_));
  XOR2_X1   g141(.A(G127gat), .B(G155gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G183gat), .B(G211gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n341_), .A2(new_n342_), .A3(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(KEYINPUT17), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n341_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n327_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n291_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355_));
  INV_X1    g154(.A(G183gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT25), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(G183gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT26), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n360_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G169gat), .ZN(new_n367_));
  INV_X1    g166(.A(G176gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(KEYINPUT79), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(G169gat), .B2(G176gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n369_), .A2(new_n371_), .A3(KEYINPUT24), .A4(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n355_), .B1(new_n366_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT78), .B(G190gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n364_), .B1(new_n376_), .B2(KEYINPUT26), .ZN(new_n377_));
  OAI211_X1 g176(.A(KEYINPUT80), .B(new_n373_), .C1(new_n377_), .C2(new_n360_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(G183gat), .B2(G190gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(G183gat), .A3(G190gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT81), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n383_), .A2(new_n379_), .A3(G183gat), .A4(G190gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT24), .B1(new_n369_), .B2(new_n371_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n375_), .A2(new_n378_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G190gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT23), .B1(new_n356_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n381_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(G183gat), .B2(new_n376_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(G169gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n388_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT84), .B(G204gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G197gat), .ZN(new_n398_));
  INV_X1    g197(.A(G197gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT83), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G197gat), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n400_), .A2(new_n402_), .A3(KEYINPUT86), .A4(G204gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n398_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT83), .B(G197gat), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT86), .B1(new_n405_), .B2(G204gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G211gat), .B(G218gat), .Z(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT21), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT21), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n407_), .B2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(G204gat), .B1(new_n400_), .B2(new_n402_), .ZN(new_n413_));
  INV_X1    g212(.A(G204gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT84), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G204gat), .ZN(new_n417_));
  AOI21_X1  g216(.A(G197gat), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT21), .B1(new_n413_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT85), .B(KEYINPUT21), .C1(new_n413_), .C2(new_n418_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n410_), .B1(new_n412_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT91), .B1(new_n396_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n405_), .A2(G204gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n428_), .A2(new_n411_), .A3(new_n398_), .A4(new_n403_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n408_), .ZN(new_n430_));
  OAI22_X1  g229(.A1(G197gat), .A2(new_n397_), .B1(new_n405_), .B2(G204gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT85), .B1(new_n431_), .B2(KEYINPUT21), .ZN(new_n432_));
  INV_X1    g231(.A(new_n422_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n429_), .B(new_n430_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n407_), .A2(new_n409_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT91), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n388_), .A2(new_n395_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n425_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT19), .ZN(new_n443_));
  NAND2_X1  g242(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n365_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n365_), .A2(KEYINPUT87), .A3(new_n444_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n360_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n450_));
  AND2_X1   g249(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n451_));
  AOI211_X1 g250(.A(new_n450_), .B(new_n451_), .C1(new_n369_), .C2(new_n371_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n369_), .A2(new_n371_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n372_), .B1(new_n451_), .B2(new_n450_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n391_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n449_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(G183gat), .A2(G190gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n394_), .B1(new_n385_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT89), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT89), .B(new_n394_), .C1(new_n385_), .C2(new_n457_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n456_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AOI211_X1 g261(.A(new_n441_), .B(new_n443_), .C1(new_n462_), .C2(new_n424_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n440_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n443_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n441_), .B1(new_n396_), .B2(new_n424_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(new_n461_), .ZN(new_n467_));
  OR3_X1    g266(.A1(new_n449_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n436_), .A2(new_n469_), .ZN(new_n470_));
  AOI211_X1 g269(.A(KEYINPUT90), .B(new_n465_), .C1(new_n466_), .C2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n434_), .A2(new_n435_), .A3(new_n395_), .A4(new_n388_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n473_), .B(KEYINPUT20), .C1(new_n424_), .C2(new_n462_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n474_), .B2(new_n443_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n464_), .B1(new_n471_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G8gat), .B(G36gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT18), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G64gat), .B(G92gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n464_), .B(new_n480_), .C1(new_n471_), .C2(new_n475_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT27), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n466_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n468_), .A2(new_n458_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT20), .B1(new_n436_), .B2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n425_), .B2(new_n439_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n485_), .B1(new_n488_), .B2(new_n465_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n481_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n490_), .A2(new_n483_), .A3(KEYINPUT27), .ZN(new_n491_));
  INV_X1    g290(.A(G134gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G127gat), .ZN(new_n493_));
  INV_X1    g292(.A(G127gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G134gat), .ZN(new_n495_));
  INV_X1    g294(.A(G120gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G113gat), .ZN(new_n497_));
  INV_X1    g296(.A(G113gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G120gat), .ZN(new_n499_));
  AND4_X1   g298(.A1(new_n493_), .A2(new_n495_), .A3(new_n497_), .A4(new_n499_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n493_), .A2(new_n495_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G71gat), .B(G99gat), .ZN(new_n503_));
  INV_X1    g302(.A(G43gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n388_), .A2(new_n395_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n388_), .B2(new_n395_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n502_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G227gat), .A2(G233gat), .ZN(new_n511_));
  INV_X1    g310(.A(G15gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT30), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT31), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n438_), .A2(new_n505_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n493_), .A2(new_n495_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n497_), .A2(new_n499_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n493_), .A2(new_n495_), .A3(new_n497_), .A4(new_n499_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n521_), .A3(new_n507_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n510_), .A2(new_n515_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n515_), .B1(new_n510_), .B2(new_n522_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G155gat), .A2(G162gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G155gat), .A2(G162gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n529_), .B1(new_n533_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(G141gat), .ZN(new_n539_));
  INV_X1    g338(.A(G148gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G141gat), .A2(G148gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n526_), .B1(KEYINPUT1), .B2(new_n528_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT1), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(G155gat), .A3(G162gat), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n538_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT3), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT2), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n542_), .A2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n553_), .A2(new_n555_), .A3(new_n534_), .A4(new_n530_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n528_), .A3(new_n527_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n528_), .A2(KEYINPUT1), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n527_), .A2(new_n558_), .A3(new_n546_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT28), .B1(new_n561_), .B2(KEYINPUT29), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n551_), .A2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n436_), .B(new_n563_), .C1(new_n550_), .C2(new_n548_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n548_), .A2(new_n550_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n562_), .B(new_n551_), .C1(new_n424_), .C2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(G233gat), .ZN(new_n567_));
  INV_X1    g366(.A(G228gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT82), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT82), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(G228gat), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n567_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(G78gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(G106gat), .ZN(new_n574_));
  INV_X1    g373(.A(G78gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n572_), .B(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n226_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G22gat), .B(G50gat), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n574_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n564_), .A2(new_n566_), .A3(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n584_));
  OAI22_X1  g383(.A1(new_n524_), .A2(new_n525_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n510_), .A2(new_n522_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n515_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n564_), .A2(new_n566_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n582_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n564_), .A2(new_n566_), .A3(new_n582_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n588_), .A2(new_n591_), .A3(new_n592_), .A4(new_n523_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n585_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n502_), .B1(new_n538_), .B2(new_n547_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT94), .B(KEYINPUT4), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n557_), .A2(new_n521_), .A3(new_n560_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(KEYINPUT4), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n595_), .A2(new_n598_), .A3(KEYINPUT92), .A4(KEYINPUT4), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n597_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G225gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT93), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n595_), .A2(new_n598_), .A3(new_n604_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G57gat), .B(G85gat), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G1gat), .B(G29gat), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n614_), .A2(new_n615_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n611_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n610_), .A3(new_n616_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n609_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n606_), .A2(new_n608_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n594_), .A2(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n484_), .A2(new_n491_), .A3(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n583_), .A2(new_n584_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n524_), .A2(new_n525_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n464_), .B(new_n635_), .C1(new_n471_), .C2(new_n475_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n473_), .A2(KEYINPUT20), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n462_), .A2(new_n424_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n443_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT90), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n474_), .A2(new_n472_), .A3(new_n443_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n644_), .A2(KEYINPUT98), .A3(new_n464_), .A4(new_n635_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n635_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n489_), .A2(new_n646_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n638_), .A2(new_n645_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n607_), .B(new_n622_), .C1(new_n603_), .C2(new_n605_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(KEYINPUT97), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT97), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n625_), .A2(new_n652_), .A3(KEYINPUT33), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n603_), .A2(new_n604_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n595_), .A2(new_n598_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n605_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n655_), .B(new_n622_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n482_), .A2(new_n654_), .A3(new_n483_), .A4(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n634_), .B1(new_n648_), .B2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n629_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n336_), .A2(new_n337_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n304_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(G229gat), .A2(G233gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n338_), .A2(new_n301_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n338_), .A2(new_n301_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(new_n665_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT77), .B(new_n666_), .C1(new_n668_), .C2(new_n664_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(KEYINPUT77), .B2(new_n666_), .ZN(new_n670_));
  XOR2_X1   g469(.A(G113gat), .B(G141gat), .Z(new_n671_));
  XNOR2_X1  g470(.A(G169gat), .B(G197gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n670_), .B(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n661_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n354_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT99), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n678_), .A2(KEYINPUT99), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n627_), .A2(G1gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT38), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n680_), .A2(KEYINPUT38), .A3(new_n679_), .A4(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n648_), .A2(new_n659_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n633_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n490_), .A2(new_n483_), .A3(KEYINPUT27), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n626_), .B1(new_n585_), .B2(new_n593_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n482_), .A2(new_n483_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n688_), .B(new_n689_), .C1(new_n690_), .C2(KEYINPUT27), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n687_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n319_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT100), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n285_), .A2(new_n675_), .A3(new_n351_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G1gat), .B1(new_n696_), .B2(new_n627_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n684_), .A2(new_n685_), .A3(new_n697_), .ZN(G1324gat));
  NOR2_X1   g497(.A1(new_n484_), .A2(new_n491_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(G8gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n680_), .A2(new_n679_), .A3(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G8gat), .B1(new_n696_), .B2(new_n699_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(KEYINPUT39), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(KEYINPUT39), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n701_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT40), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n701_), .B(KEYINPUT40), .C1(new_n703_), .C2(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1325gat));
  INV_X1    g508(.A(new_n632_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G15gat), .B1(new_n696_), .B2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT41), .Z(new_n712_));
  NAND3_X1  g511(.A1(new_n678_), .A2(new_n512_), .A3(new_n632_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1326gat));
  OR3_X1    g513(.A1(new_n677_), .A2(G22gat), .A3(new_n630_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G22gat), .B1(new_n696_), .B2(new_n630_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n716_), .A2(KEYINPUT42), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(KEYINPUT42), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n715_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT101), .Z(G1327gat));
  INV_X1    g519(.A(new_n351_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(new_n319_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n676_), .A2(new_n284_), .A3(new_n722_), .ZN(new_n723_));
  OR3_X1    g522(.A1(new_n723_), .A2(G29gat), .A3(new_n627_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n284_), .A2(new_n674_), .A3(new_n351_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n284_), .A2(KEYINPUT102), .A3(new_n674_), .A4(new_n351_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n692_), .B2(new_n327_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n731_), .B(new_n327_), .C1(new_n629_), .C2(new_n660_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n725_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n327_), .B1(new_n629_), .B2(new_n660_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT43), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n739_), .A2(new_n733_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n627_), .B1(new_n737_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n735_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n740_), .A2(KEYINPUT103), .ZN(new_n747_));
  AND4_X1   g546(.A1(new_n744_), .A2(new_n746_), .A3(new_n747_), .A4(new_n736_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT44), .B1(new_n735_), .B2(new_n745_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n744_), .B1(new_n749_), .B2(new_n747_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n742_), .B(new_n743_), .C1(new_n748_), .C2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G29gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n747_), .A3(new_n736_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT104), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n749_), .A2(new_n744_), .A3(new_n747_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n743_), .B1(new_n756_), .B2(new_n742_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n724_), .B1(new_n752_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(G1328gat));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n761_));
  INV_X1    g560(.A(new_n723_), .ZN(new_n762_));
  INV_X1    g561(.A(G36gat), .ZN(new_n763_));
  INV_X1    g562(.A(new_n699_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n699_), .B1(new_n737_), .B2(new_n741_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n769_), .B2(G36gat), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT109), .B(new_n761_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773_));
  INV_X1    g572(.A(new_n767_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n735_), .A2(new_n725_), .A3(new_n736_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT105), .B1(new_n740_), .B2(KEYINPUT44), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n764_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n778_), .B2(new_n763_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n773_), .B1(new_n779_), .B2(KEYINPUT108), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT46), .B1(new_n770_), .B2(KEYINPUT109), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n772_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(G1329gat));
  NOR2_X1   g582(.A1(new_n775_), .A2(new_n776_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n784_), .A2(new_n504_), .A3(new_n710_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n756_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(KEYINPUT110), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n762_), .A2(new_n632_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT110), .B1(new_n788_), .B2(new_n504_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n785_), .B2(new_n756_), .ZN(new_n790_));
  XOR2_X1   g589(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n791_));
  OR3_X1    g590(.A1(new_n787_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1330gat));
  AOI211_X1 g593(.A(new_n630_), .B(new_n784_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n795_));
  INV_X1    g594(.A(G50gat), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n630_), .A2(G50gat), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT112), .ZN(new_n798_));
  OAI22_X1  g597(.A1(new_n795_), .A2(new_n796_), .B1(new_n723_), .B2(new_n798_), .ZN(G1331gat));
  NOR2_X1   g598(.A1(new_n661_), .A2(new_n674_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n800_), .A2(new_n285_), .A3(new_n352_), .ZN(new_n801_));
  AOI21_X1  g600(.A(G57gat), .B1(new_n801_), .B2(new_n626_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n674_), .A2(new_n351_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n694_), .A2(new_n290_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n233_), .B1(new_n626_), .B2(KEYINPUT113), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(KEYINPUT113), .B2(new_n233_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n802_), .B1(new_n804_), .B2(new_n806_), .ZN(G1332gat));
  AOI21_X1  g606(.A(new_n231_), .B1(new_n804_), .B2(new_n764_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n801_), .A2(new_n231_), .A3(new_n764_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1333gat));
  INV_X1    g611(.A(G71gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n804_), .B2(new_n632_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n801_), .A2(new_n813_), .A3(new_n632_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(G1334gat));
  AOI21_X1  g617(.A(new_n575_), .B1(new_n804_), .B2(new_n631_), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n819_), .B(KEYINPUT50), .Z(new_n820_));
  NAND3_X1  g619(.A1(new_n801_), .A2(new_n575_), .A3(new_n631_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1335gat));
  NAND3_X1  g621(.A1(new_n290_), .A2(new_n722_), .A3(new_n800_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n823_), .A2(G85gat), .A3(new_n627_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n285_), .A2(new_n675_), .A3(new_n351_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n739_), .B2(new_n733_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n626_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n824_), .B1(G85gat), .B2(new_n827_), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT116), .Z(G1336gat));
  INV_X1    g628(.A(new_n823_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G92gat), .B1(new_n830_), .B2(new_n764_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n764_), .A2(new_n221_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n826_), .B2(new_n832_), .ZN(G1337gat));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT51), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n632_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n823_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(G99gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n826_), .B2(new_n632_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n840_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n837_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n834_), .A2(KEYINPUT51), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1338gat));
  AOI21_X1  g644(.A(new_n226_), .B1(new_n826_), .B2(new_n631_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT52), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n823_), .A2(G106gat), .A3(new_n630_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(KEYINPUT53), .Z(G1339gat));
  XNOR2_X1  g649(.A(new_n803_), .B(KEYINPUT119), .ZN(new_n851_));
  INV_X1    g650(.A(new_n327_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n284_), .A3(new_n852_), .ZN(new_n853_));
  XOR2_X1   g652(.A(new_n853_), .B(KEYINPUT54), .Z(new_n854_));
  INV_X1    g653(.A(new_n319_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n259_), .A2(new_n207_), .A3(new_n262_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n276_), .A2(KEYINPUT55), .A3(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(new_n205_), .C1(KEYINPUT55), .C2(new_n276_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT56), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n859_), .ZN(new_n861_));
  OR3_X1    g660(.A1(new_n860_), .A2(new_n861_), .A3(KEYINPUT120), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n860_), .B2(KEYINPUT120), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n279_), .A2(new_n280_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n674_), .A4(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n281_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n663_), .A2(new_n665_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n664_), .B1(new_n867_), .B2(KEYINPUT121), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(KEYINPUT121), .B2(new_n867_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n668_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n673_), .B1(new_n870_), .B2(new_n664_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n670_), .A2(new_n673_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n866_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n855_), .B1(new_n865_), .B2(new_n873_), .ZN(new_n874_));
  OR3_X1    g673(.A1(new_n874_), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n864_), .B(new_n872_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n852_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n874_), .A2(KEYINPUT57), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT122), .B1(new_n874_), .B2(KEYINPUT57), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n875_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n854_), .B1(new_n882_), .B2(new_n351_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n764_), .A2(new_n627_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n593_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n883_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G113gat), .B1(new_n888_), .B2(new_n674_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n874_), .A2(KEYINPUT57), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n721_), .B1(new_n890_), .B2(new_n880_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n891_), .A2(new_n854_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n887_), .A2(KEYINPUT59), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n888_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n674_), .A2(G113gat), .ZN(new_n898_));
  XOR2_X1   g697(.A(new_n898_), .B(KEYINPUT123), .Z(new_n899_));
  AOI21_X1  g698(.A(new_n889_), .B1(new_n897_), .B2(new_n899_), .ZN(G1340gat));
  OAI21_X1  g699(.A(G120gat), .B1(new_n896_), .B2(new_n291_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n883_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n886_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n904_));
  AOI21_X1  g703(.A(G120gat), .B1(new_n285_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT124), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n904_), .B2(G120gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n905_), .B2(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n901_), .B1(new_n903_), .B2(new_n909_), .ZN(G1341gat));
  AOI21_X1  g709(.A(G127gat), .B1(new_n888_), .B2(new_n721_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n494_), .B1(new_n721_), .B2(KEYINPUT125), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(KEYINPUT125), .B2(new_n494_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n897_), .B2(new_n913_), .ZN(G1342gat));
  NOR3_X1   g713(.A1(new_n883_), .A2(new_n319_), .A3(new_n887_), .ZN(new_n915_));
  OAI21_X1  g714(.A(KEYINPUT126), .B1(new_n915_), .B2(G134gat), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n917_), .B(new_n492_), .C1(new_n903_), .C2(new_n319_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n852_), .A2(new_n492_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n916_), .A2(new_n918_), .B1(new_n897_), .B2(new_n919_), .ZN(G1343gat));
  NOR2_X1   g719(.A1(new_n883_), .A2(new_n585_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n674_), .A3(new_n884_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g722(.A1(new_n921_), .A2(new_n290_), .A3(new_n884_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g724(.A1(new_n921_), .A2(new_n721_), .A3(new_n884_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT61), .B(G155gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1346gat));
  INV_X1    g727(.A(G162gat), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n921_), .A2(new_n929_), .A3(new_n855_), .A4(new_n884_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n921_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n931_), .A2(new_n852_), .A3(new_n885_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n930_), .B1(new_n932_), .B2(new_n929_), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n699_), .A2(new_n626_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n593_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n892_), .A2(new_n674_), .A3(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT62), .B1(new_n937_), .B2(KEYINPUT22), .ZN(new_n938_));
  OAI21_X1  g737(.A(G169gat), .B1(new_n937_), .B2(KEYINPUT62), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n940_), .B1(new_n367_), .B2(new_n938_), .ZN(G1348gat));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n883_), .A2(new_n593_), .A3(new_n935_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n291_), .A2(new_n368_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n942_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n892_), .A2(new_n936_), .ZN(new_n946_));
  AOI21_X1  g745(.A(G176gat), .B1(new_n946_), .B2(new_n285_), .ZN(new_n947_));
  AND4_X1   g746(.A1(new_n942_), .A2(new_n902_), .A3(new_n936_), .A4(new_n944_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n945_), .A2(new_n947_), .A3(new_n948_), .ZN(G1349gat));
  AOI21_X1  g748(.A(G183gat), .B1(new_n943_), .B2(new_n721_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n351_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n946_), .B2(new_n951_), .ZN(G1350gat));
  AOI21_X1  g751(.A(new_n319_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n946_), .A2(new_n953_), .ZN(new_n954_));
  AND2_X1   g753(.A1(new_n946_), .A2(new_n327_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n955_), .B2(new_n389_), .ZN(G1351gat));
  NAND3_X1  g755(.A1(new_n921_), .A2(new_n674_), .A3(new_n934_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g757(.A1(new_n921_), .A2(new_n290_), .A3(new_n934_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n959_), .A2(new_n397_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n960_), .B1(new_n414_), .B2(new_n959_), .ZN(G1353gat));
  XOR2_X1   g760(.A(KEYINPUT63), .B(G211gat), .Z(new_n962_));
  AND4_X1   g761(.A1(new_n721_), .A2(new_n921_), .A3(new_n934_), .A4(new_n962_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n921_), .A2(new_n721_), .A3(new_n934_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n963_), .B1(new_n964_), .B2(new_n965_), .ZN(G1354gat));
  INV_X1    g765(.A(G218gat), .ZN(new_n967_));
  NAND4_X1  g766(.A1(new_n921_), .A2(new_n967_), .A3(new_n855_), .A4(new_n934_), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n931_), .A2(new_n852_), .A3(new_n935_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n968_), .B1(new_n969_), .B2(new_n967_), .ZN(G1355gat));
endmodule


