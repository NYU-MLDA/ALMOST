//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n929_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_, new_n976_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G197gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(G197gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT21), .B1(new_n204_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT83), .B1(new_n203_), .B2(G204gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT83), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(new_n205_), .A3(G197gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n209_), .B(new_n211_), .C1(G197gat), .C2(new_n205_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n207_), .B(new_n208_), .C1(new_n212_), .C2(KEYINPUT21), .ZN(new_n213_));
  INV_X1    g012(.A(new_n208_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(KEYINPUT21), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT82), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G155gat), .B(G162gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT3), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(KEYINPUT2), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(KEYINPUT2), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n217_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n220_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(KEYINPUT1), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(G155gat), .A3(G162gat), .ZN(new_n230_));
  AOI211_X1 g029(.A(new_n218_), .B(new_n225_), .C1(new_n228_), .C2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT29), .B1(new_n224_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n202_), .B1(new_n216_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n216_), .A2(new_n232_), .A3(new_n202_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G78gat), .B(G106gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT85), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n240_));
  NOR2_X1   g039(.A1(new_n224_), .A2(new_n231_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT29), .ZN(new_n242_));
  XOR2_X1   g041(.A(G22gat), .B(G50gat), .Z(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n240_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n246_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n240_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n244_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n216_), .A2(new_n232_), .A3(new_n202_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n236_), .B1(new_n252_), .B2(new_n233_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT85), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n234_), .A2(new_n254_), .A3(new_n235_), .A4(new_n237_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n239_), .A2(new_n251_), .A3(new_n253_), .A4(new_n255_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n252_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT84), .B(new_n236_), .C1(new_n252_), .C2(new_n233_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n257_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n256_), .B1(new_n261_), .B2(new_n251_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT86), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n256_), .B(KEYINPUT86), .C1(new_n261_), .C2(new_n251_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G113gat), .B(G120gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT79), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n269_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G113gat), .B(G120gat), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n268_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT79), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n218_), .A2(KEYINPUT3), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n218_), .A2(KEYINPUT3), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n279_), .A2(new_n280_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n228_), .A2(new_n230_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n225_), .A2(new_n218_), .ZN(new_n283_));
  OAI22_X1  g082(.A1(new_n281_), .A2(new_n217_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n272_), .A2(new_n278_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT93), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n274_), .A2(new_n276_), .A3(new_n271_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n271_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n291_), .A2(KEYINPUT93), .A3(new_n285_), .A4(new_n284_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n272_), .A2(new_n278_), .A3(new_n284_), .A4(KEYINPUT91), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n241_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT91), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(new_n241_), .B2(new_n270_), .ZN(new_n297_));
  OAI211_X1 g096(.A(KEYINPUT4), .B(new_n294_), .C1(new_n295_), .C2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G225gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT92), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n293_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G29gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n303_), .B(KEYINPUT0), .Z(new_n304_));
  INV_X1    g103(.A(G57gat), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n305_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n306_), .A2(G85gat), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(G85gat), .B1(new_n306_), .B2(new_n307_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n291_), .A2(new_n284_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT91), .B1(new_n284_), .B2(new_n277_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n300_), .A3(new_n294_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n302_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G8gat), .B(G36gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G64gat), .B(G92gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT25), .B(G183gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT88), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT26), .B(G190gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(KEYINPUT24), .A3(new_n332_), .ZN(new_n333_));
  OR3_X1    g132(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(G183gat), .A4(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT23), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(G183gat), .A3(G190gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(KEYINPUT76), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n335_), .A2(new_n338_), .A3(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT89), .ZN(new_n346_));
  INV_X1    g145(.A(new_n332_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G169gat), .ZN(new_n348_));
  INV_X1    g147(.A(G176gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n345_), .A2(KEYINPUT89), .ZN(new_n352_));
  OAI22_X1  g151(.A1(new_n330_), .A2(new_n343_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n213_), .A2(new_n215_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n325_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n354_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n342_), .A2(new_n338_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n350_), .B1(new_n357_), .B2(new_n344_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n340_), .A2(new_n341_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n328_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G190gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n360_), .B1(new_n362_), .B2(KEYINPUT26), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n326_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n335_), .B(new_n359_), .C1(new_n361_), .C2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n356_), .A2(new_n358_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n324_), .B1(new_n355_), .B2(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n335_), .A2(new_n338_), .A3(new_n342_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT88), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n326_), .B(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n328_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n351_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n352_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n356_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n365_), .A2(new_n358_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n354_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n324_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(new_n325_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n321_), .B1(new_n367_), .B2(new_n382_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n371_), .A2(new_n368_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n366_), .B(KEYINPUT20), .C1(new_n384_), .C2(new_n356_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n379_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n320_), .A3(new_n381_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n315_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT33), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT95), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n301_), .B(new_n294_), .C1(new_n295_), .C2(new_n297_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT94), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n313_), .A2(KEYINPUT94), .A3(new_n301_), .A4(new_n294_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n301_), .B1(new_n288_), .B2(new_n292_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n394_), .A2(new_n395_), .B1(new_n396_), .B2(new_n298_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n310_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n391_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n395_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n298_), .ZN(new_n401_));
  AND4_X1   g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n398_), .A4(new_n391_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n388_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n401_), .A3(new_n398_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n397_), .A2(new_n398_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n320_), .A2(KEYINPUT32), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n386_), .A2(new_n381_), .A3(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n377_), .B2(new_n354_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n324_), .B1(new_n411_), .B2(new_n376_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n356_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n377_), .A2(new_n354_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n325_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n412_), .B1(new_n415_), .B2(new_n324_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n409_), .B1(new_n416_), .B2(new_n408_), .ZN(new_n417_));
  OAI22_X1  g216(.A1(new_n403_), .A2(KEYINPUT96), .B1(new_n407_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n315_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n404_), .A2(new_n390_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n397_), .A2(new_n398_), .A3(new_n391_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT96), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n267_), .B1(new_n418_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n291_), .B(KEYINPUT31), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n377_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G15gat), .B(G43gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT77), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G71gat), .B(G99gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n431_), .B(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n365_), .A2(new_n358_), .A3(KEYINPUT30), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n428_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT78), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n428_), .A2(new_n435_), .A3(KEYINPUT78), .A4(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n428_), .A2(new_n436_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n435_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n426_), .B1(new_n445_), .B2(KEYINPUT80), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT80), .ZN(new_n447_));
  INV_X1    g246(.A(new_n426_), .ZN(new_n448_));
  AOI211_X1 g247(.A(new_n447_), .B(new_n448_), .C1(new_n441_), .C2(new_n444_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n264_), .A2(new_n450_), .A3(new_n265_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n425_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT98), .B1(new_n405_), .B2(new_n406_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n400_), .A2(new_n401_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n310_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT98), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n404_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n387_), .A2(KEYINPUT27), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n416_), .A2(new_n320_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n383_), .A2(new_n387_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT27), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  OAI22_X1  g266(.A1(new_n451_), .A2(new_n452_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n454_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT65), .ZN(new_n470_));
  OAI22_X1  g269(.A1(new_n470_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(KEYINPUT7), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n470_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(KEYINPUT8), .A3(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n483_));
  INV_X1    g282(.A(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(KEYINPUT9), .A3(new_n480_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n480_), .A2(KEYINPUT9), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n476_), .A2(new_n486_), .A3(new_n487_), .A4(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n482_), .A2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT8), .B1(new_n478_), .B2(new_n481_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G57gat), .B(G64gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G71gat), .B(G78gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(KEYINPUT11), .ZN(new_n495_));
  INV_X1    g294(.A(G64gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G57gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n305_), .A2(G64gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n498_), .A3(KEYINPUT11), .ZN(new_n499_));
  AND2_X1   g298(.A1(G71gat), .A2(G78gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G71gat), .A2(G78gat), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n495_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n492_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n499_), .A2(new_n502_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n503_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G230gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT64), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT12), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n514_), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT12), .B(new_n510_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n517_), .A2(new_n506_), .A3(new_n518_), .A4(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G120gat), .B(G148gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT5), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G176gat), .B(G204gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n525_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n515_), .A2(new_n520_), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT66), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(KEYINPUT13), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(KEYINPUT13), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n526_), .A2(new_n530_), .A3(KEYINPUT13), .A4(new_n528_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(G1gat), .ZN(new_n541_));
  INV_X1    g340(.A(G8gat), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT14), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(G22gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(G15gat), .ZN(new_n545_));
  INV_X1    g344(.A(G15gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(G22gat), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(KEYINPUT71), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G1gat), .B(G8gat), .Z(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(KEYINPUT71), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n551_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n552_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n554_), .B1(new_n555_), .B2(new_n549_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G29gat), .B(G36gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT68), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G43gat), .B(G50gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT73), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n557_), .A2(KEYINPUT68), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(KEYINPUT68), .ZN(new_n563_));
  INV_X1    g362(.A(new_n559_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n560_), .A2(new_n561_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n561_), .B1(new_n560_), .B2(new_n565_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n553_), .B(new_n556_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n560_), .A2(new_n565_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT73), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n556_), .A2(new_n553_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n560_), .A2(new_n561_), .A3(new_n565_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n568_), .A2(new_n570_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n565_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n564_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT15), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT15), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n560_), .A2(new_n580_), .A3(new_n565_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n556_), .A2(new_n553_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n570_), .B1(new_n584_), .B2(new_n575_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n540_), .B1(new_n576_), .B2(new_n585_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n573_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n569_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n568_), .A2(new_n570_), .A3(new_n575_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n539_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(KEYINPUT74), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT74), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n589_), .A2(new_n593_), .A3(new_n590_), .A4(new_n539_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n469_), .A2(new_n536_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n505_), .B(new_n597_), .Z(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n573_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n505_), .B(new_n597_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n583_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G127gat), .B(G155gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT16), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n599_), .A2(new_n601_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT72), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n599_), .A2(new_n607_), .A3(new_n601_), .A4(KEYINPUT72), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n605_), .B(KEYINPUT17), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n599_), .A2(new_n601_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT36), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT35), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n490_), .A2(new_n491_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n582_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT69), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n625_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n492_), .A2(new_n571_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n624_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT35), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n627_), .A2(new_n630_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n629_), .A2(new_n634_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n582_), .A2(new_n626_), .B1(new_n632_), .B2(new_n631_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT69), .B1(new_n582_), .B2(new_n626_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n636_), .B(new_n630_), .C1(new_n637_), .C2(new_n625_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n621_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT70), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n620_), .A2(KEYINPUT36), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n639_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n642_), .ZN(new_n644_));
  AOI221_X4 g443(.A(new_n640_), .B1(new_n644_), .B2(new_n621_), .C1(new_n635_), .C2(new_n638_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT37), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n639_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n635_), .A2(new_n638_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT70), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n649_), .A3(new_n644_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n641_), .B1(new_n639_), .B2(new_n642_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n646_), .A2(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n596_), .A2(new_n616_), .A3(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n541_), .A3(new_n460_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT38), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n643_), .A2(new_n645_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n469_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n595_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n661_), .A2(new_n535_), .A3(new_n616_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n460_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n657_), .A2(new_n665_), .ZN(G1324gat));
  NAND3_X1  g465(.A1(new_n660_), .A2(new_n467_), .A3(new_n662_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G8gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT99), .B1(new_n668_), .B2(KEYINPUT39), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n667_), .A2(new_n670_), .A3(new_n671_), .A4(G8gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n668_), .A2(KEYINPUT39), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n669_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n655_), .A2(new_n542_), .A3(new_n467_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n674_), .A2(KEYINPUT40), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1325gat));
  INV_X1    g479(.A(new_n450_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G15gat), .B1(new_n663_), .B2(new_n681_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n683_));
  OR2_X1    g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n683_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n655_), .A2(new_n546_), .A3(new_n450_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n684_), .A2(new_n685_), .A3(new_n686_), .ZN(G1326gat));
  OAI21_X1  g486(.A(G22gat), .B1(new_n663_), .B2(new_n267_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n655_), .A2(new_n544_), .A3(new_n266_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1327gat));
  INV_X1    g491(.A(new_n596_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n616_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n658_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n664_), .A2(G29gat), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT106), .Z(new_n697_));
  NAND3_X1  g496(.A1(new_n693_), .A2(new_n695_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n661_), .A2(new_n535_), .A3(new_n694_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT102), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n417_), .B1(new_n457_), .B2(new_n404_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n403_), .A2(KEYINPUT96), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n266_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n266_), .A2(new_n681_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n264_), .A2(new_n450_), .A3(new_n265_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n468_), .B(new_n654_), .C1(new_n705_), .C2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(KEYINPUT43), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n454_), .A2(new_n712_), .A3(new_n468_), .A4(new_n654_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n710_), .B1(new_n709_), .B2(KEYINPUT43), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n701_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT44), .B(new_n701_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n460_), .A4(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(G29gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n718_), .A2(new_n460_), .A3(new_n720_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT104), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n699_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  AND4_X1   g524(.A1(new_n699_), .A2(new_n724_), .A3(G29gat), .A4(new_n721_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n698_), .B1(new_n725_), .B2(new_n726_), .ZN(G1328gat));
  NAND2_X1  g526(.A1(new_n693_), .A2(new_n695_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n467_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(G36gat), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n718_), .A2(new_n467_), .A3(new_n720_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G36gat), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(KEYINPUT46), .A3(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1329gat));
  NOR3_X1   g539(.A1(new_n728_), .A2(G43gat), .A3(new_n681_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n718_), .A2(new_n450_), .A3(new_n720_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G43gat), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g543(.A1(new_n718_), .A2(G50gat), .A3(new_n266_), .A4(new_n720_), .ZN(new_n745_));
  INV_X1    g544(.A(G50gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n728_), .B2(new_n267_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1331gat));
  AOI21_X1  g547(.A(new_n616_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n660_), .A2(new_n535_), .A3(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G57gat), .B1(new_n750_), .B2(new_n664_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n536_), .A2(new_n595_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n469_), .A2(new_n752_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n753_), .A2(new_n616_), .A3(new_n654_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n305_), .A3(new_n460_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n751_), .A2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT107), .ZN(G1332gat));
  OAI21_X1  g556(.A(G64gat), .B1(new_n750_), .B2(new_n729_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT48), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n754_), .A2(new_n496_), .A3(new_n467_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n750_), .B2(new_n681_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT49), .ZN(new_n763_));
  INV_X1    g562(.A(G71gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n754_), .A2(new_n764_), .A3(new_n450_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1334gat));
  OAI21_X1  g565(.A(G78gat), .B1(new_n750_), .B2(new_n267_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n754_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n267_), .A2(G78gat), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT109), .Z(new_n772_));
  OAI21_X1  g571(.A(new_n769_), .B1(new_n770_), .B2(new_n772_), .ZN(G1335gat));
  OR2_X1    g572(.A1(new_n714_), .A2(new_n715_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n752_), .A2(new_n616_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT110), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(G85gat), .B1(new_n777_), .B2(new_n664_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n753_), .A2(new_n658_), .A3(new_n694_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n664_), .A2(G85gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n780_), .B2(new_n781_), .ZN(G1336gat));
  AOI21_X1  g581(.A(G92gat), .B1(new_n779_), .B2(new_n467_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n777_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n467_), .A2(G92gat), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT111), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n784_), .B2(new_n786_), .ZN(G1337gat));
  NAND4_X1  g586(.A1(new_n779_), .A2(new_n450_), .A3(new_n483_), .A4(new_n485_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n774_), .A2(new_n450_), .A3(new_n776_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n789_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT112), .B1(new_n789_), .B2(G99gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n788_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT51), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n788_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n779_), .A2(new_n484_), .A3(new_n266_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n774_), .A2(new_n266_), .A3(new_n776_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT53), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(new_n797_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1339gat));
  NAND2_X1  g605(.A1(new_n729_), .A2(new_n460_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT119), .B1(new_n807_), .B2(new_n707_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n807_), .A2(KEYINPUT119), .A3(new_n707_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n810_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n808_), .A3(KEYINPUT120), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT59), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  XOR2_X1   g615(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n817_));
  NAND3_X1  g616(.A1(new_n584_), .A2(new_n570_), .A3(new_n575_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n568_), .A2(new_n575_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n539_), .B(new_n818_), .C1(new_n819_), .C2(new_n570_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n586_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n529_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n528_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n490_), .A2(new_n510_), .A3(new_n491_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n516_), .B2(new_n511_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n827_), .B2(new_n519_), .ZN(new_n828_));
  AND4_X1   g627(.A1(new_n825_), .A2(new_n517_), .A3(new_n506_), .A4(new_n519_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n514_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n520_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n520_), .A2(new_n835_), .A3(new_n831_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n520_), .B2(new_n831_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n525_), .B1(new_n834_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n517_), .A2(new_n506_), .A3(new_n519_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT116), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n517_), .A2(new_n506_), .A3(new_n825_), .A4(new_n519_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n832_), .B1(new_n845_), .B2(new_n514_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n520_), .A2(new_n831_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT115), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n520_), .A2(new_n835_), .A3(new_n831_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(KEYINPUT56), .A3(new_n525_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n824_), .B1(new_n841_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n823_), .B1(new_n853_), .B2(new_n595_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n658_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n817_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT56), .B1(new_n851_), .B2(new_n525_), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n840_), .B(new_n527_), .C1(new_n846_), .C2(new_n850_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n528_), .B(new_n595_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n822_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(KEYINPUT57), .A3(new_n658_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n856_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n528_), .B(new_n821_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT58), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n841_), .A2(new_n852_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n528_), .A4(new_n821_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n654_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n694_), .B1(new_n862_), .B2(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n643_), .A2(KEYINPUT37), .A3(new_n645_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n651_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n749_), .A2(new_n534_), .A3(new_n533_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n873_), .A2(KEYINPUT113), .A3(new_n874_), .A4(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n875_), .A2(new_n646_), .A3(new_n874_), .A4(new_n653_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT113), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n536_), .A2(new_n749_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n654_), .B2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n876_), .A2(new_n879_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n876_), .A2(new_n879_), .A3(KEYINPUT114), .A4(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n816_), .B1(new_n870_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n595_), .A2(G113gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT121), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n873_), .B1(new_n864_), .B2(new_n867_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n856_), .B(new_n861_), .C1(KEYINPUT118), .C2(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n890_), .A2(KEYINPUT118), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n616_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n884_), .A2(new_n885_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n811_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n887_), .B(new_n889_), .C1(new_n895_), .C2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(G113gat), .B1(new_n895_), .B2(new_n595_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1340gat));
  OAI211_X1 g699(.A(new_n535_), .B(new_n887_), .C1(new_n895_), .C2(new_n896_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G120gat), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n903_));
  INV_X1    g702(.A(G120gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n535_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n895_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n902_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT122), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n902_), .A2(new_n910_), .A3(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1341gat));
  OAI21_X1  g711(.A(new_n887_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT124), .B(G127gat), .ZN(new_n914_));
  OR3_X1    g713(.A1(new_n913_), .A2(new_n616_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(G127gat), .B1(new_n895_), .B2(new_n694_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n916_), .A2(new_n917_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n915_), .A2(new_n918_), .A3(new_n919_), .ZN(G1342gat));
  OAI21_X1  g719(.A(G134gat), .B1(new_n913_), .B2(new_n873_), .ZN(new_n921_));
  INV_X1    g720(.A(G134gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n895_), .A2(new_n922_), .A3(new_n855_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1343gat));
  AND2_X1   g723(.A1(new_n893_), .A2(new_n894_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n925_), .A2(new_n706_), .A3(new_n807_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n595_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n535_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g729(.A1(new_n926_), .A2(new_n694_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT61), .B(G155gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1346gat));
  INV_X1    g732(.A(G162gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n926_), .A2(new_n934_), .A3(new_n855_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n926_), .A2(new_n654_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n934_), .ZN(G1347gat));
  AND2_X1   g736(.A1(new_n862_), .A2(new_n869_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n894_), .B1(new_n938_), .B2(new_n694_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n664_), .A2(new_n467_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n681_), .ZN(new_n941_));
  XOR2_X1   g740(.A(new_n941_), .B(KEYINPUT125), .Z(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n266_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n939_), .A2(new_n943_), .ZN(new_n944_));
  OAI21_X1  g743(.A(G169gat), .B1(new_n944_), .B2(new_n661_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n945_), .A2(KEYINPUT62), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(KEYINPUT62), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n595_), .A2(new_n348_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(KEYINPUT126), .ZN(new_n949_));
  OAI22_X1  g748(.A1(new_n946_), .A2(new_n947_), .B1(new_n944_), .B2(new_n949_), .ZN(G1348gat));
  NOR2_X1   g749(.A1(new_n925_), .A2(new_n266_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n942_), .A2(new_n349_), .A3(new_n536_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n939_), .A2(new_n535_), .A3(new_n943_), .ZN(new_n953_));
  AOI22_X1  g752(.A1(new_n951_), .A2(new_n952_), .B1(new_n953_), .B2(new_n349_), .ZN(G1349gat));
  NOR2_X1   g753(.A1(new_n942_), .A2(new_n616_), .ZN(new_n955_));
  AOI21_X1  g754(.A(G183gat), .B1(new_n951_), .B2(new_n955_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n944_), .A2(new_n370_), .A3(new_n616_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1350gat));
  OAI21_X1  g757(.A(G190gat), .B1(new_n944_), .B2(new_n873_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n855_), .A2(new_n328_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n944_), .B2(new_n960_), .ZN(G1351gat));
  NOR3_X1   g760(.A1(new_n925_), .A2(new_n706_), .A3(new_n940_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(new_n595_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n535_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n967_));
  INV_X1    g766(.A(G211gat), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n694_), .B1(new_n967_), .B2(new_n968_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(KEYINPUT127), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n962_), .A2(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n967_), .A2(new_n968_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n971_), .B(new_n972_), .ZN(G1354gat));
  INV_X1    g772(.A(G218gat), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n962_), .A2(new_n974_), .A3(new_n855_), .ZN(new_n975_));
  AND2_X1   g774(.A1(new_n962_), .A2(new_n654_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n975_), .B1(new_n976_), .B2(new_n974_), .ZN(G1355gat));
endmodule


