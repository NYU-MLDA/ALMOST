//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT84), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n210_), .B(new_n211_), .C1(G183gat), .C2(G190gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n202_), .A2(KEYINPUT84), .A3(new_n203_), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n206_), .A2(new_n207_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT83), .ZN(new_n216_));
  INV_X1    g015(.A(G190gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(KEYINPUT26), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n215_), .B(new_n218_), .C1(new_n219_), .C2(new_n216_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n208_), .B(new_n209_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n203_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(KEYINPUT24), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n220_), .A2(new_n222_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G211gat), .B(G218gat), .Z(new_n228_));
  INV_X1    g027(.A(KEYINPUT21), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n230_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n228_), .A3(KEYINPUT21), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n214_), .A2(new_n227_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT20), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT95), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT95), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n239_), .A3(KEYINPUT20), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n234_), .A2(new_n235_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n224_), .A2(new_n207_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n215_), .A2(new_n219_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n223_), .A3(new_n203_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n245_), .A2(new_n222_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT97), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n202_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT22), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(G169gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n223_), .A2(KEYINPUT22), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT97), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n255_), .A3(new_n203_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n207_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT98), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT99), .B1(new_n221_), .B2(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n212_), .A2(KEYINPUT99), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n257_), .A2(new_n258_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n256_), .A2(KEYINPUT98), .A3(new_n207_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n249_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n238_), .B(new_n240_), .C1(new_n242_), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G8gat), .B(G36gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n214_), .A2(new_n227_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n241_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n267_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n276_), .A2(KEYINPUT20), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n257_), .A2(new_n258_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n261_), .A2(new_n260_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n263_), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(new_n242_), .A3(new_n248_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n268_), .A2(new_n274_), .A3(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n284_), .A2(KEYINPUT27), .ZN(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT104), .B(KEYINPUT20), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n288_), .A2(KEYINPUT105), .B1(new_n241_), .B2(new_n275_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n286_), .B1(new_n264_), .B2(new_n242_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT105), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n277_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n265_), .A2(new_n267_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n273_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n236_), .A2(new_n239_), .A3(KEYINPUT20), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n239_), .B1(new_n236_), .B2(KEYINPUT20), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n281_), .A2(new_n248_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n241_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n277_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n283_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n273_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n284_), .ZN(new_n304_));
  XOR2_X1   g103(.A(KEYINPUT106), .B(KEYINPUT27), .Z(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n285_), .A2(new_n295_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT102), .B(KEYINPUT0), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT103), .ZN(new_n309_));
  XOR2_X1   g108(.A(G1gat), .B(G29gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G57gat), .B(G85gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316_));
  INV_X1    g115(.A(G141gat), .ZN(new_n317_));
  INV_X1    g116(.A(G148gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G155gat), .B(G162gat), .Z(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(KEYINPUT89), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT89), .B1(new_n324_), .B2(new_n325_), .ZN(new_n328_));
  INV_X1    g127(.A(G155gat), .ZN(new_n329_));
  INV_X1    g128(.A(G162gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT1), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G155gat), .A3(G162gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n330_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G141gat), .B(G148gat), .Z(new_n336_));
  AND3_X1   g135(.A1(new_n335_), .A2(KEYINPUT88), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT88), .B1(new_n335_), .B2(new_n336_), .ZN(new_n338_));
  OAI22_X1  g137(.A1(new_n327_), .A2(new_n328_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G127gat), .B(G134gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT86), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n341_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G113gat), .B(G120gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n339_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n324_), .A2(new_n325_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n326_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n335_), .A2(new_n336_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT88), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n335_), .A2(KEYINPUT88), .A3(new_n336_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n354_), .A2(new_n359_), .A3(new_n348_), .A4(new_n347_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n350_), .A2(new_n360_), .A3(KEYINPUT4), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n354_), .A2(new_n359_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT101), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AND4_X1   g163(.A1(KEYINPUT101), .A2(new_n339_), .A3(new_n349_), .A4(new_n363_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n315_), .B(new_n361_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n350_), .A2(new_n360_), .A3(new_n314_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n313_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n366_), .A2(new_n367_), .A3(new_n313_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n353_), .A2(new_n326_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n241_), .B(new_n373_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n242_), .B1(new_n339_), .B2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n378_), .B2(new_n373_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n380_), .B(KEYINPUT93), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n376_), .B(new_n381_), .C1(new_n378_), .C2(new_n373_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT91), .ZN(new_n386_));
  XOR2_X1   g185(.A(G22gat), .B(G50gat), .Z(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n339_), .B2(KEYINPUT29), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n374_), .A2(new_n375_), .A3(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n386_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n391_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n339_), .A2(KEYINPUT29), .A3(new_n387_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n389_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(KEYINPUT91), .A3(new_n392_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n395_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n392_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n402_), .A2(new_n384_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT94), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n379_), .A2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n376_), .B(KEYINPUT94), .C1(new_n378_), .C2(new_n373_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n380_), .A3(new_n406_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n385_), .A2(new_n401_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409_));
  INV_X1    g208(.A(G71gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G99gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n275_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(new_n349_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G15gat), .B(G43gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT85), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT30), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n417_), .B(KEYINPUT31), .Z(new_n418_));
  XNOR2_X1  g217(.A(new_n414_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n307_), .A2(new_n372_), .A3(new_n408_), .A4(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n370_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n314_), .B(new_n361_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n313_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n350_), .A2(new_n360_), .A3(new_n315_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n423_), .A2(new_n303_), .A3(new_n284_), .A4(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n370_), .A2(new_n422_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n274_), .A2(KEYINPUT32), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n268_), .A2(new_n283_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n370_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(new_n368_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n276_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n288_), .A2(KEYINPUT105), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n267_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n294_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n430_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n428_), .A2(new_n429_), .B1(new_n433_), .B2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n408_), .A2(new_n371_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n439_), .A2(new_n408_), .B1(new_n307_), .B2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n419_), .B(KEYINPUT87), .Z(new_n442_));
  OAI21_X1  g241(.A(new_n421_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G29gat), .B(G36gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT74), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G43gat), .B(G50gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT78), .B(G8gat), .ZN(new_n448_));
  INV_X1    g247(.A(G1gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT14), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G15gat), .B(G22gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G1gat), .B(G8gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT80), .B1(new_n447_), .B2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n447_), .A2(new_n457_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(G229gat), .A3(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n447_), .B(KEYINPUT15), .ZN(new_n462_));
  INV_X1    g261(.A(new_n457_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n447_), .A2(new_n457_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G229gat), .A2(G233gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT81), .Z(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n461_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G113gat), .B(G141gat), .Z(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT82), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G169gat), .B(G197gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n461_), .A2(new_n468_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n443_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G230gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G99gat), .A2(G106gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT6), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(G99gat), .A3(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT66), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(G99gat), .ZN(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT67), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT7), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n492_), .A2(new_n488_), .A3(new_n489_), .A4(KEYINPUT67), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n482_), .A2(new_n484_), .A3(KEYINPUT66), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n487_), .A2(new_n491_), .A3(new_n493_), .A4(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G85gat), .B(G92gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(KEYINPUT8), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n491_), .A2(new_n485_), .A3(new_n493_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n496_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT8), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(G85gat), .A3(G92gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(new_n496_), .B2(new_n504_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT65), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT65), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n508_), .B(new_n505_), .C1(new_n496_), .C2(new_n504_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n511_));
  OR2_X1    g310(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n487_), .A2(new_n494_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n503_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G64gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(G57gat), .ZN(new_n520_));
  INV_X1    g319(.A(G57gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(G64gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT68), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT11), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT70), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n521_), .A2(G64gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n519_), .A2(G57gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT68), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(KEYINPUT11), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n527_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT11), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n536_), .A3(new_n531_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT69), .ZN(new_n538_));
  XOR2_X1   g337(.A(G71gat), .B(G78gat), .Z(new_n539_));
  AND3_X1   g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n535_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT69), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n544_), .A2(new_n545_), .B1(new_n527_), .B2(new_n534_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n518_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n544_), .A2(new_n527_), .A3(new_n534_), .A4(new_n545_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n533_), .B1(new_n532_), .B2(KEYINPUT11), .ZN(new_n549_));
  AOI211_X1 g348(.A(KEYINPUT70), .B(new_n536_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n550_));
  OAI22_X1  g349(.A1(new_n540_), .A2(new_n541_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n498_), .A2(new_n502_), .B1(new_n510_), .B2(new_n516_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(KEYINPUT12), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n552_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n480_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n548_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(new_n555_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(new_n479_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(G176gat), .B(G204gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT72), .ZN(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n562_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT13), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n572_), .A2(KEYINPUT13), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT73), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(KEYINPUT73), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n457_), .B(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n548_), .A2(new_n551_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G127gat), .B(G155gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589_));
  OR3_X1    g388(.A1(new_n588_), .A2(KEYINPUT79), .A3(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n584_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n589_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n584_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n462_), .A2(new_n518_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT34), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT35), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n552_), .A2(new_n447_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n596_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n599_), .A2(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n604_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n596_), .A2(new_n606_), .A3(new_n601_), .A4(new_n602_), .ZN(new_n607_));
  XOR2_X1   g406(.A(G190gat), .B(G218gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT75), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT77), .Z(new_n614_));
  AND3_X1   g413(.A1(new_n605_), .A2(new_n607_), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n611_), .B(KEYINPUT36), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n615_), .A2(new_n617_), .A3(KEYINPUT37), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT37), .B1(new_n615_), .B2(new_n617_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AND4_X1   g420(.A1(new_n478_), .A2(new_n580_), .A3(new_n595_), .A4(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n449_), .A3(new_n371_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT38), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n615_), .A2(new_n617_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n443_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n576_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n477_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n627_), .A2(new_n594_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n449_), .B1(new_n630_), .B2(new_n371_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n625_), .A2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(new_n624_), .B2(new_n623_), .ZN(G1324gat));
  INV_X1    g432(.A(new_n307_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n622_), .A2(new_n634_), .A3(new_n448_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n630_), .A2(new_n634_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n636_), .A2(new_n637_), .A3(G8gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n636_), .B2(G8gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(G1325gat));
  INV_X1    g441(.A(G15gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n630_), .B2(new_n442_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT107), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT107), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT41), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT41), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n622_), .A2(new_n643_), .A3(new_n442_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT108), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n649_), .A3(new_n651_), .ZN(G1326gat));
  INV_X1    g451(.A(G22gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n408_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n622_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n630_), .B2(new_n654_), .ZN(new_n656_));
  XOR2_X1   g455(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(G1327gat));
  INV_X1    g459(.A(new_n626_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n594_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n576_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n478_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G29gat), .B1(new_n665_), .B2(new_n371_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n629_), .A2(new_n595_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n443_), .A2(new_n668_), .A3(new_n620_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n443_), .B2(new_n620_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n667_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT44), .B(new_n667_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n371_), .A2(G29gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n666_), .B1(new_n675_), .B2(new_n676_), .ZN(G1328gat));
  NOR2_X1   g476(.A1(new_n307_), .A2(G36gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n478_), .A2(new_n663_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n478_), .A2(KEYINPUT45), .A3(new_n663_), .A4(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n673_), .A2(new_n634_), .A3(new_n674_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(G36gat), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(KEYINPUT110), .A3(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(KEYINPUT110), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n686_), .A2(KEYINPUT110), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n685_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n687_), .A2(new_n690_), .ZN(G1329gat));
  NAND4_X1  g490(.A1(new_n673_), .A2(G43gat), .A3(new_n420_), .A4(new_n674_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n442_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n664_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(G43gat), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g495(.A(G50gat), .B1(new_n665_), .B2(new_n654_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n654_), .A2(G50gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n675_), .B2(new_n698_), .ZN(G1331gat));
  INV_X1    g498(.A(new_n627_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n477_), .A2(new_n594_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n700_), .A2(new_n579_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G57gat), .B1(new_n703_), .B2(new_n372_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n477_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n443_), .A2(new_n705_), .ZN(new_n706_));
  AND4_X1   g505(.A1(new_n576_), .A2(new_n706_), .A3(new_n595_), .A4(new_n621_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(new_n521_), .A3(new_n371_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n704_), .A2(new_n708_), .ZN(G1332gat));
  NAND3_X1  g508(.A1(new_n707_), .A2(new_n519_), .A3(new_n634_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n702_), .A2(new_n634_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(G64gat), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n711_), .B2(G64gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT112), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n717_), .B(new_n710_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1333gat));
  NAND3_X1  g518(.A1(new_n707_), .A2(new_n410_), .A3(new_n442_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT49), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n702_), .A2(new_n442_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(G71gat), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT49), .B(new_n410_), .C1(new_n702_), .C2(new_n442_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT113), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(new_n720_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1334gat));
  INV_X1    g528(.A(G78gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n702_), .B2(new_n654_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT50), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n707_), .A2(new_n730_), .A3(new_n654_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1335gat));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n580_), .A2(new_n662_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(new_n706_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n662_), .ZN(new_n739_));
  AND4_X1   g538(.A1(new_n735_), .A2(new_n706_), .A3(new_n579_), .A4(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G85gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n743_), .A3(new_n371_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n576_), .A2(new_n705_), .A3(new_n594_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n670_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n443_), .A2(new_n668_), .A3(new_n620_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(KEYINPUT115), .A3(new_n747_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n745_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(KEYINPUT116), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n754_), .B(new_n745_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n753_), .A2(new_n755_), .A3(new_n372_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n744_), .B1(new_n756_), .B2(new_n743_), .ZN(G1336gat));
  INV_X1    g556(.A(G92gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n742_), .A2(new_n758_), .A3(new_n634_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n753_), .A2(new_n755_), .A3(new_n307_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n758_), .ZN(G1337gat));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n511_), .A2(new_n513_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n420_), .B(new_n763_), .C1(new_n737_), .C2(new_n740_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n752_), .A2(new_n442_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n762_), .B(new_n764_), .C1(new_n765_), .C2(new_n488_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n764_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n488_), .B1(new_n752_), .B2(new_n442_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT51), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(G1338gat));
  AND3_X1   g569(.A1(new_n654_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n737_), .B2(new_n740_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n745_), .A2(new_n408_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n748_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n489_), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n774_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n772_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n772_), .B(new_n781_), .C1(new_n778_), .C2(new_n777_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n621_), .A2(new_n701_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n576_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n628_), .A2(KEYINPUT118), .A3(new_n621_), .A4(new_n701_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(KEYINPUT54), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n784_), .B(new_n789_), .C1(new_n785_), .C2(new_n576_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n460_), .A2(new_n467_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n467_), .B1(new_n447_), .B2(new_n457_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n475_), .B1(new_n464_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n476_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n571_), .B2(new_n569_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n554_), .A2(new_n557_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT55), .A3(new_n479_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n558_), .A2(KEYINPUT120), .A3(KEYINPUT55), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  AOI211_X1 g604(.A(KEYINPUT12), .B(new_n552_), .C1(new_n548_), .C2(new_n551_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n560_), .B2(KEYINPUT12), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT119), .B(new_n805_), .C1(new_n807_), .C2(new_n480_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n558_), .B2(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n807_), .A2(new_n480_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n804_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n570_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n568_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n799_), .A2(new_n479_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT119), .B1(new_n819_), .B2(new_n805_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n558_), .A2(new_n809_), .A3(KEYINPUT55), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n812_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n803_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT120), .B1(new_n558_), .B2(KEYINPUT55), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n818_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT122), .ZN(new_n827_));
  INV_X1    g626(.A(new_n818_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n808_), .A2(new_n810_), .B1(new_n480_), .B2(new_n807_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n804_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n816_), .A2(new_n827_), .A3(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n477_), .A2(new_n569_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n798_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n792_), .B1(new_n835_), .B2(new_n661_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n568_), .B1(new_n829_), .B2(new_n804_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n815_), .ZN(new_n838_));
  OAI22_X1  g637(.A1(new_n831_), .A2(new_n830_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n826_), .A2(KEYINPUT122), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n834_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n798_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n626_), .A2(KEYINPUT57), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n797_), .B1(new_n562_), .B2(new_n568_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n570_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT58), .B(new_n847_), .C1(new_n848_), .C2(new_n830_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n620_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n851_));
  OAI21_X1  g650(.A(new_n826_), .B1(new_n837_), .B2(KEYINPUT56), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n847_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n850_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n836_), .A2(new_n846_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n791_), .B1(new_n855_), .B2(new_n594_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n634_), .A2(new_n654_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(new_n371_), .A3(new_n420_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(G113gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n477_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT57), .B1(new_n843_), .B2(new_n626_), .ZN(new_n864_));
  OAI22_X1  g663(.A1(new_n835_), .A2(new_n844_), .B1(new_n853_), .B2(new_n850_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n594_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n791_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n858_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(KEYINPUT59), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n705_), .B1(new_n863_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n861_), .B1(new_n871_), .B2(new_n860_), .ZN(G1340gat));
  INV_X1    g671(.A(G120gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n628_), .B2(KEYINPUT60), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n859_), .B(new_n874_), .C1(KEYINPUT60), .C2(new_n873_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n580_), .B1(new_n863_), .B2(new_n870_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n873_), .ZN(G1341gat));
  INV_X1    g676(.A(G127gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n859_), .A2(new_n878_), .A3(new_n595_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n594_), .B1(new_n863_), .B2(new_n870_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n878_), .ZN(G1342gat));
  INV_X1    g680(.A(G134gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n859_), .A2(new_n882_), .A3(new_n661_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n621_), .B1(new_n863_), .B2(new_n870_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n882_), .ZN(G1343gat));
  NOR2_X1   g684(.A1(new_n442_), .A2(new_n408_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n887_), .A2(new_n634_), .A3(new_n372_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n868_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n317_), .A3(new_n477_), .ZN(new_n891_));
  OAI21_X1  g690(.A(G141gat), .B1(new_n889_), .B2(new_n705_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1344gat));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n318_), .A3(new_n579_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G148gat), .B1(new_n889_), .B2(new_n580_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1345gat));
  NAND3_X1  g695(.A1(new_n868_), .A2(new_n595_), .A3(new_n888_), .ZN(new_n897_));
  XOR2_X1   g696(.A(KEYINPUT61), .B(G155gat), .Z(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT124), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n897_), .B(new_n899_), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n889_), .B2(new_n621_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n661_), .A2(new_n330_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n889_), .B2(new_n902_), .ZN(G1347gat));
  AND3_X1   g702(.A1(new_n477_), .A2(new_n255_), .A3(new_n251_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n307_), .A2(new_n371_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n907_), .A2(new_n693_), .A3(new_n654_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n868_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n908_), .ZN(new_n910_));
  AOI211_X1 g709(.A(KEYINPUT126), .B(new_n910_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n904_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n913_));
  AOI211_X1 g712(.A(new_n705_), .B(new_n910_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n223_), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n913_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n913_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n868_), .A2(new_n908_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n915_), .B(new_n918_), .C1(new_n919_), .C2(new_n705_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n912_), .A2(new_n917_), .A3(new_n920_), .ZN(G1348gat));
  OAI211_X1 g720(.A(new_n203_), .B(new_n576_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n922_));
  OAI21_X1  g721(.A(G176gat), .B1(new_n919_), .B2(new_n580_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1349gat));
  NOR2_X1   g723(.A1(new_n856_), .A2(new_n910_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G183gat), .B1(new_n925_), .B2(new_n595_), .ZN(new_n926_));
  OAI21_X1  g725(.A(KEYINPUT126), .B1(new_n856_), .B2(new_n910_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n868_), .A2(new_n905_), .A3(new_n908_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n594_), .A2(new_n215_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n926_), .B1(new_n929_), .B2(new_n930_), .ZN(G1350gat));
  AND2_X1   g730(.A1(new_n661_), .A2(new_n219_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n932_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n621_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n934_), .B2(new_n217_), .ZN(G1351gat));
  NOR2_X1   g734(.A1(new_n887_), .A2(new_n907_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n856_), .A2(new_n937_), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n938_), .A2(G197gat), .A3(new_n477_), .ZN(new_n939_));
  AOI21_X1  g738(.A(G197gat), .B1(new_n938_), .B2(new_n477_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1352gat));
  NAND2_X1  g740(.A1(new_n868_), .A2(new_n936_), .ZN(new_n942_));
  OAI211_X1 g741(.A(KEYINPUT127), .B(G204gat), .C1(new_n942_), .C2(new_n580_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n938_), .A2(new_n579_), .A3(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n945_), .ZN(G1353gat));
  OR2_X1    g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n947_), .B1(new_n938_), .B2(new_n595_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n942_), .A2(new_n594_), .ZN(new_n949_));
  XOR2_X1   g748(.A(KEYINPUT63), .B(G211gat), .Z(new_n950_));
  AOI21_X1  g749(.A(new_n948_), .B1(new_n949_), .B2(new_n950_), .ZN(G1354gat));
  OR3_X1    g750(.A1(new_n942_), .A2(G218gat), .A3(new_n626_), .ZN(new_n952_));
  OAI21_X1  g751(.A(G218gat), .B1(new_n942_), .B2(new_n621_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1355gat));
endmodule


