//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G64gat), .B(G92gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT91), .ZN(new_n212_));
  INV_X1    g011(.A(G197gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n212_), .B1(new_n213_), .B2(G204gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n211_), .A2(KEYINPUT21), .A3(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G197gat), .B(G204gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n211_), .A2(KEYINPUT21), .ZN(new_n218_));
  XOR2_X1   g017(.A(G197gat), .B(G204gat), .Z(new_n219_));
  NAND4_X1  g018(.A1(new_n219_), .A2(KEYINPUT21), .A3(new_n211_), .A4(new_n214_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G183gat), .ZN(new_n222_));
  INV_X1    g021(.A(G190gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT23), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT81), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n223_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT81), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n229_), .B(KEYINPUT23), .C1(new_n222_), .C2(new_n223_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  INV_X1    g032(.A(G176gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n232_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G183gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n222_), .A2(KEYINPUT25), .ZN(new_n239_));
  AND2_X1   g038(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n238_), .B(new_n239_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT94), .ZN(new_n243_));
  INV_X1    g042(.A(G169gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n234_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(KEYINPUT24), .A3(new_n232_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(new_n243_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT83), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n248_), .B(KEYINPUT23), .C1(new_n222_), .C2(new_n223_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT83), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n245_), .A2(KEYINPUT24), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n247_), .A2(new_n249_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n243_), .B1(new_n242_), .B2(new_n246_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n221_), .B(new_n236_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT20), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n227_), .A2(new_n230_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n238_), .A2(KEYINPUT80), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n240_), .A2(new_n241_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n238_), .A2(new_n239_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n257_), .B(new_n258_), .C1(new_n259_), .C2(KEYINPUT80), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n256_), .A2(new_n260_), .A3(new_n251_), .A4(new_n246_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n250_), .A2(new_n228_), .A3(new_n249_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT82), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n235_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n233_), .A2(KEYINPUT82), .A3(new_n234_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n262_), .A2(new_n264_), .A3(new_n232_), .A4(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n221_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n210_), .B1(new_n255_), .B2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n236_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n221_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n261_), .A2(new_n266_), .A3(new_n221_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n271_), .A2(KEYINPUT20), .A3(new_n272_), .A4(new_n209_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n207_), .B1(new_n268_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n209_), .B1(new_n255_), .B2(new_n267_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n271_), .A2(KEYINPUT20), .A3(new_n272_), .A4(new_n210_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n207_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n279_), .A3(KEYINPUT27), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT27), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n268_), .A2(new_n273_), .A3(new_n207_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(new_n274_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G141gat), .ZN(new_n293_));
  INV_X1    g092(.A(G148gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(new_n292_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n298_));
  NOR2_X1   g097(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n291_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT89), .ZN(new_n301_));
  AND3_X1   g100(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT87), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n293_), .B(new_n294_), .C1(new_n303_), .C2(KEYINPUT3), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n305_), .B(KEYINPUT87), .C1(G141gat), .C2(G148gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT89), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n308_), .B(new_n291_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n286_), .A2(new_n288_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n297_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n270_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(G228gat), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G78gat), .B(G106gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n270_), .B(new_n318_), .C1(new_n312_), .C2(new_n322_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n320_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT93), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n320_), .A2(new_n323_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n321_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT93), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n320_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n312_), .A2(new_n322_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G22gat), .B(G50gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT28), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n333_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n326_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(KEYINPUT93), .C1(new_n324_), .C2(new_n325_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT104), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n310_), .A2(new_n311_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n296_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G127gat), .A2(G134gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(G113gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G127gat), .A2(G134gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n347_), .ZN(new_n349_));
  OAI21_X1  g148(.A(G113gat), .B1(new_n349_), .B2(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G120gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n348_), .A2(new_n350_), .A3(G120gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n343_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n312_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(KEYINPUT4), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT98), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT97), .B(KEYINPUT4), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n343_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n361_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n348_), .A2(new_n350_), .A3(G120gat), .ZN(new_n365_));
  AOI21_X1  g164(.A(G120gat), .B1(new_n348_), .B2(new_n350_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT98), .B1(new_n312_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT96), .Z(new_n371_));
  NAND3_X1  g170(.A1(new_n359_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT0), .B(G57gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G85gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(G1gat), .B(G29gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n312_), .B(new_n355_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n371_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n372_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n376_), .B1(new_n372_), .B2(new_n379_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n285_), .A2(new_n340_), .A3(new_n341_), .A4(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT104), .B1(new_n385_), .B2(new_n284_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT103), .ZN(new_n389_));
  INV_X1    g188(.A(new_n207_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(new_n268_), .B2(new_n273_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n278_), .A2(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT102), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT102), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n278_), .A2(new_n398_), .A3(new_n392_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n389_), .B1(new_n395_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n372_), .A2(new_n379_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n376_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n393_), .B1(new_n404_), .B2(new_n380_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n398_), .B1(new_n278_), .B2(new_n392_), .ZN(new_n406_));
  AOI211_X1 g205(.A(KEYINPUT102), .B(new_n391_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(KEYINPUT103), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n401_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n380_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT99), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT99), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n380_), .A2(new_n414_), .A3(new_n411_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n282_), .A2(new_n274_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n372_), .A2(KEYINPUT33), .A3(new_n376_), .A4(new_n379_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT100), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n359_), .A2(new_n369_), .A3(new_n378_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n376_), .B1(new_n377_), .B2(new_n371_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n419_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n417_), .B(new_n418_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT101), .B1(new_n416_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n415_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n414_), .B1(new_n380_), .B2(new_n411_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT101), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n410_), .B1(new_n425_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n388_), .B1(new_n432_), .B2(new_n340_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n261_), .A2(new_n266_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n434_), .A2(KEYINPUT30), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(KEYINPUT30), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n357_), .B1(new_n439_), .B2(KEYINPUT84), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n438_), .A2(new_n441_), .A3(new_n355_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n444_), .B(KEYINPUT86), .Z(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n439_), .A2(KEYINPUT84), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G71gat), .B(G99gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G15gat), .B(G43gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(G227gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n446_), .B1(new_n447_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n438_), .A2(new_n441_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n452_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n454_), .A2(new_n445_), .A3(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n443_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n447_), .A2(new_n446_), .A3(new_n452_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n445_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n442_), .A4(new_n440_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT105), .B1(new_n340_), .B2(new_n284_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n383_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT105), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n338_), .A2(new_n339_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n285_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n463_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT106), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT106), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n463_), .A2(new_n465_), .A3(new_n468_), .A4(new_n471_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n433_), .A2(new_n462_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G120gat), .B(G148gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G176gat), .B(G204gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT6), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n482_));
  OR3_X1    g281(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT8), .ZN(new_n485_));
  XOR2_X1   g284(.A(G85gat), .B(G92gat), .Z(new_n486_));
  AND3_X1   g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT10), .B(G99gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(G106gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT65), .ZN(new_n491_));
  NOR2_X1   g290(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n493_), .B1(KEYINPUT9), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G92gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n486_), .A2(KEYINPUT9), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n481_), .A3(new_n497_), .ZN(new_n498_));
  OAI22_X1  g297(.A1(new_n487_), .A2(new_n488_), .B1(new_n491_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT68), .ZN(new_n500_));
  XOR2_X1   g299(.A(G57gat), .B(G64gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT67), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G57gat), .B(G64gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n500_), .B1(new_n506_), .B2(KEYINPUT11), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT11), .ZN(new_n508_));
  AOI211_X1 g307(.A(KEYINPUT68), .B(new_n508_), .C1(new_n502_), .C2(new_n505_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n502_), .A2(new_n508_), .A3(new_n505_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G71gat), .B(G78gat), .Z(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n507_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n503_), .B(KEYINPUT67), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT68), .B1(new_n514_), .B2(new_n508_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n506_), .A2(new_n500_), .A3(KEYINPUT11), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n515_), .A2(new_n516_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n499_), .B1(new_n513_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n488_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT65), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n490_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n498_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n519_), .A2(new_n520_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n515_), .A2(new_n510_), .A3(new_n516_), .A4(new_n511_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n512_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n499_), .B2(KEYINPUT69), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n518_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n525_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n531_), .B(new_n499_), .C1(KEYINPUT69), .C2(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT64), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n518_), .A2(new_n527_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n535_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n479_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n539_), .A3(new_n479_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n541_), .A2(KEYINPUT13), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT13), .B1(new_n541_), .B2(new_n542_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(new_n244_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n213_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550_));
  XOR2_X1   g349(.A(G29gat), .B(G36gat), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT72), .B(G43gat), .ZN(new_n553_));
  INV_X1    g352(.A(G50gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n553_), .A2(new_n554_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n552_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT73), .ZN(new_n559_));
  XOR2_X1   g358(.A(KEYINPUT72), .B(G43gat), .Z(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G50gat), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(new_n551_), .A3(new_n555_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n558_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n559_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n550_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n558_), .A2(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT73), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n558_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(KEYINPUT15), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571_));
  INV_X1    g370(.A(G8gat), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G1gat), .B(G8gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n570_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n576_), .A2(new_n562_), .A3(new_n558_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT78), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n578_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n566_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n579_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n549_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n578_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n549_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(KEYINPUT79), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT79), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n591_), .B(new_n549_), .C1(new_n582_), .C2(new_n584_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n546_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n473_), .A2(new_n596_), .ZN(new_n597_));
  OR3_X1    g396(.A1(new_n499_), .A2(KEYINPUT74), .A3(new_n566_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT71), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT34), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT35), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT76), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT74), .B1(new_n570_), .B2(new_n499_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n499_), .A2(new_n566_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n598_), .B(new_n603_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT75), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(KEYINPUT75), .B(new_n598_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n601_), .A2(new_n602_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(G134gat), .ZN(new_n615_));
  INV_X1    g414(.A(G162gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n611_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n612_), .A2(new_n613_), .A3(new_n617_), .A4(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n613_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n617_), .A2(new_n613_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n611_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n621_), .B(new_n622_), .C1(new_n624_), .C2(new_n618_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n576_), .B(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(new_n531_), .ZN(new_n630_));
  XOR2_X1   g429(.A(G127gat), .B(G155gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT17), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n636_), .A2(KEYINPUT69), .A3(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n630_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(KEYINPUT17), .B2(new_n635_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n639_), .B1(new_n630_), .B2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n627_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n597_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT107), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n202_), .B1(new_n645_), .B2(new_n464_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT108), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n620_), .A2(KEYINPUT37), .A3(new_n625_), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT37), .B1(new_n620_), .B2(new_n625_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n642_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n597_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n202_), .A3(new_n464_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT38), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n647_), .A2(new_n654_), .ZN(G1324gat));
  OAI21_X1  g454(.A(G8gat), .B1(new_n644_), .B2(new_n285_), .ZN(new_n656_));
  XOR2_X1   g455(.A(KEYINPUT109), .B(KEYINPUT39), .Z(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n652_), .A2(new_n572_), .A3(new_n284_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g460(.A1(new_n645_), .A2(new_n461_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G15gat), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n462_), .A2(G15gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n651_), .B2(new_n666_), .ZN(G1326gat));
  INV_X1    g466(.A(G22gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n645_), .B2(new_n340_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT42), .Z(new_n670_));
  NAND3_X1  g469(.A1(new_n652_), .A2(new_n668_), .A3(new_n340_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1327gat));
  NAND2_X1  g471(.A1(new_n627_), .A2(new_n642_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT112), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n597_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n383_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT111), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n470_), .A2(new_n472_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n405_), .A2(KEYINPUT103), .A3(new_n408_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT103), .B1(new_n405_), .B2(new_n408_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n430_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n416_), .A2(new_n424_), .A3(KEYINPUT101), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n387_), .B1(new_n684_), .B2(new_n467_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n677_), .B(new_n678_), .C1(new_n685_), .C2(new_n461_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n648_), .A2(new_n649_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(KEYINPUT111), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n686_), .B(new_n688_), .C1(new_n473_), .C2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n689_), .A2(KEYINPUT110), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n689_), .A2(KEYINPUT110), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(new_n473_), .B2(new_n687_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n642_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n596_), .A2(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n691_), .A2(new_n693_), .A3(new_n695_), .A4(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n678_), .B1(new_n685_), .B2(new_n461_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n688_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n692_), .B1(new_n702_), .B2(new_n694_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n703_), .A2(KEYINPUT44), .A3(new_n691_), .A4(new_n697_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n700_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n464_), .ZN(new_n706_));
  MUX2_X1   g505(.A(new_n676_), .B(new_n706_), .S(G29gat), .Z(G1328gat));
  NOR3_X1   g506(.A1(new_n675_), .A2(G36gat), .A3(new_n285_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT45), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n700_), .A2(new_n284_), .A3(new_n704_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n710_), .A2(KEYINPUT113), .A3(G36gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT113), .B1(new_n710_), .B2(G36gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT46), .B(new_n709_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND3_X1  g516(.A1(new_n705_), .A2(G43gat), .A3(new_n461_), .ZN(new_n718_));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n675_), .B2(new_n462_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g521(.A1(new_n705_), .A2(G50gat), .A3(new_n340_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n554_), .B1(new_n675_), .B2(new_n467_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1331gat));
  NAND2_X1  g524(.A1(new_n546_), .A2(new_n594_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n473_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n650_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n464_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(new_n643_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(new_n383_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(G57gat), .B2(new_n732_), .ZN(G1332gat));
  OAI21_X1  g532(.A(G64gat), .B1(new_n731_), .B2(new_n285_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n285_), .A2(G64gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n728_), .B2(new_n736_), .ZN(G1333gat));
  OR3_X1    g536(.A1(new_n728_), .A2(G71gat), .A3(new_n462_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G71gat), .B1(new_n731_), .B2(new_n462_), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n739_), .A2(KEYINPUT114), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(KEYINPUT114), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(KEYINPUT49), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT49), .B1(new_n740_), .B2(new_n741_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n738_), .B1(new_n742_), .B2(new_n743_), .ZN(G1334gat));
  OR3_X1    g543(.A1(new_n728_), .A2(G78gat), .A3(new_n467_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G78gat), .B1(new_n731_), .B2(new_n467_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT115), .Z(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(KEYINPUT50), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(KEYINPUT50), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n726_), .A2(new_n696_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n691_), .A2(new_n693_), .A3(new_n695_), .A4(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT117), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n703_), .A2(KEYINPUT117), .A3(new_n691_), .A4(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(KEYINPUT118), .A3(new_n755_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n383_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(G85gat), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n674_), .A2(new_n727_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n383_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT116), .Z(new_n765_));
  NAND2_X1  g564(.A1(new_n761_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT119), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n761_), .A2(KEYINPUT119), .A3(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1336gat));
  AND3_X1   g569(.A1(new_n758_), .A2(new_n284_), .A3(new_n759_), .ZN(new_n771_));
  INV_X1    g570(.A(G92gat), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n284_), .A2(new_n772_), .ZN(new_n773_));
  OAI22_X1  g572(.A1(new_n771_), .A2(new_n772_), .B1(new_n763_), .B2(new_n773_), .ZN(G1337gat));
  OR3_X1    g573(.A1(new_n763_), .A2(new_n489_), .A3(new_n462_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n754_), .A2(new_n461_), .A3(new_n755_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT120), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G99gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G99gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT51), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n782_), .B(new_n775_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1338gat));
  OR3_X1    g583(.A1(new_n763_), .A2(G106gat), .A3(new_n467_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n752_), .A2(new_n467_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(G106gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G106gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT53), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n785_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1339gat));
  NOR2_X1   g593(.A1(new_n533_), .A2(new_n536_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n537_), .A2(KEYINPUT55), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n533_), .A2(new_n797_), .A3(new_n536_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n795_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n479_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n797_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n801_));
  AOI211_X1 g600(.A(KEYINPUT55), .B(new_n535_), .C1(new_n530_), .C2(new_n532_), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n801_), .A2(new_n802_), .B1(new_n536_), .B2(new_n533_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n478_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n593_), .A2(new_n800_), .A3(new_n542_), .A4(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n581_), .A2(new_n583_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n579_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n578_), .A2(new_n581_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n808_), .B(new_n549_), .C1(new_n579_), .C2(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n810_), .A2(new_n589_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n542_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n540_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n806_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n626_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n479_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n804_), .B1(new_n803_), .B2(new_n478_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(KEYINPUT58), .A3(new_n542_), .A4(new_n811_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n800_), .A2(new_n542_), .A3(new_n811_), .A4(new_n805_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n821_), .B(new_n824_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n814_), .A2(KEYINPUT57), .A3(new_n626_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n817_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n642_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n650_), .A2(new_n829_), .A3(new_n594_), .A4(new_n545_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT37), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n626_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n620_), .A2(KEYINPUT37), .A3(new_n625_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n594_), .A3(new_n696_), .A4(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT54), .B1(new_n834_), .B2(new_n546_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n830_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n828_), .A2(new_n836_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n463_), .A2(new_n461_), .A3(new_n468_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n464_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n383_), .B1(new_n828_), .B2(new_n836_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(KEYINPUT59), .A3(new_n838_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n845_), .A2(new_n346_), .A3(new_n594_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n346_), .B1(new_n839_), .B2(new_n594_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(KEYINPUT121), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n847_), .A2(KEYINPUT121), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n846_), .A2(new_n848_), .A3(new_n849_), .ZN(G1340gat));
  AOI21_X1  g649(.A(KEYINPUT122), .B1(new_n844_), .B2(new_n546_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n852_), .B(new_n545_), .C1(new_n841_), .C2(new_n843_), .ZN(new_n853_));
  OAI21_X1  g652(.A(G120gat), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n839_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT60), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n545_), .B2(G120gat), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n855_), .B(new_n857_), .C1(new_n856_), .C2(G120gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n858_), .ZN(G1341gat));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  AND4_X1   g659(.A1(KEYINPUT59), .A2(new_n837_), .A3(new_n464_), .A4(new_n838_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT59), .B1(new_n842_), .B2(new_n838_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n696_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G127gat), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n839_), .A2(G127gat), .A3(new_n642_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n860_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n867_));
  AOI211_X1 g666(.A(KEYINPUT123), .B(new_n865_), .C1(new_n863_), .C2(G127gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1342gat));
  AOI21_X1  g668(.A(G134gat), .B1(new_n855_), .B2(new_n627_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n845_), .A2(new_n687_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(G134gat), .ZN(G1343gat));
  AOI211_X1 g671(.A(new_n461_), .B(new_n467_), .C1(new_n828_), .C2(new_n836_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n284_), .A2(new_n383_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n594_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT124), .B(G141gat), .Z(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1344gat));
  NOR2_X1   g677(.A1(new_n875_), .A2(new_n545_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n294_), .ZN(G1345gat));
  NOR2_X1   g679(.A1(new_n875_), .A2(new_n642_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT125), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n881_), .B(new_n883_), .ZN(G1346gat));
  NOR3_X1   g683(.A1(new_n875_), .A2(new_n616_), .A3(new_n687_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n873_), .A2(new_n627_), .A3(new_n874_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n616_), .B2(new_n886_), .ZN(G1347gat));
  AND2_X1   g686(.A1(new_n837_), .A2(new_n465_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n285_), .A2(new_n340_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n593_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G169gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT126), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n893_), .A3(G169gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(KEYINPUT62), .A3(new_n894_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n888_), .A2(new_n593_), .A3(new_n233_), .A4(new_n889_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n891_), .A2(KEYINPUT126), .A3(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(new_n896_), .A3(new_n898_), .ZN(G1348gat));
  NAND2_X1  g698(.A1(new_n888_), .A2(new_n889_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n545_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n234_), .ZN(G1349gat));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n642_), .ZN(new_n903_));
  MUX2_X1   g702(.A(G183gat), .B(new_n259_), .S(new_n903_), .Z(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n900_), .B2(new_n687_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n627_), .A2(new_n258_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT127), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n900_), .B2(new_n907_), .ZN(G1351gat));
  AOI211_X1 g707(.A(new_n461_), .B(new_n385_), .C1(new_n828_), .C2(new_n836_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n284_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n594_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n213_), .ZN(G1352gat));
  INV_X1    g711(.A(new_n910_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n546_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g714(.A1(new_n910_), .A2(new_n642_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n916_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n917_));
  XOR2_X1   g716(.A(KEYINPUT63), .B(G211gat), .Z(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n916_), .B2(new_n918_), .ZN(G1354gat));
  AOI21_X1  g718(.A(G218gat), .B1(new_n913_), .B2(new_n627_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n910_), .A2(new_n687_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(G218gat), .B2(new_n921_), .ZN(G1355gat));
endmodule


