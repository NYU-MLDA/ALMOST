//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n972_, new_n973_, new_n975_, new_n976_, new_n977_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n990_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n997_, new_n998_, new_n999_;
  AND3_X1   g000(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n202_));
  AOI21_X1  g001(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209_));
  INV_X1    g008(.A(G176gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(new_n214_), .ZN(new_n215_));
  OR3_X1    g014(.A1(new_n206_), .A2(KEYINPUT76), .A3(KEYINPUT26), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT26), .B1(new_n206_), .B2(KEYINPUT76), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n212_), .A2(new_n210_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT24), .A3(new_n222_), .ZN(new_n223_));
  OR3_X1    g022(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n204_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n215_), .B1(new_n220_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G71gat), .B(G99gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(G43gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n226_), .B(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G127gat), .B(G134gat), .Z(new_n230_));
  XOR2_X1   g029(.A(G113gat), .B(G120gat), .Z(new_n231_));
  XOR2_X1   g030(.A(new_n230_), .B(new_n231_), .Z(new_n232_));
  XNOR2_X1  g031(.A(new_n229_), .B(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G227gat), .A2(G233gat), .ZN(new_n234_));
  INV_X1    g033(.A(G15gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT30), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT31), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n233_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G141gat), .A2(G148gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT2), .ZN(new_n244_));
  NAND3_X1  g043(.A1(KEYINPUT77), .A2(G141gat), .A3(G148gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n247_));
  INV_X1    g046(.A(G141gat), .ZN(new_n248_));
  INV_X1    g047(.A(G148gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT3), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n247_), .A2(new_n252_), .A3(new_n248_), .A4(new_n249_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n246_), .A2(new_n251_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G155gat), .A2(G162gat), .ZN(new_n256_));
  OR2_X1    g055(.A1(G155gat), .A2(G162gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n248_), .A2(new_n249_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n243_), .A2(new_n245_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT78), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n256_), .A2(new_n261_), .A3(KEYINPUT1), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n262_), .B(new_n257_), .C1(KEYINPUT1), .C2(new_n256_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n256_), .B2(KEYINPUT1), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n259_), .B(new_n260_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n258_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT86), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n258_), .A2(KEYINPUT80), .A3(new_n265_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .A4(new_n232_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n258_), .A2(KEYINPUT80), .A3(new_n265_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT80), .B1(new_n258_), .B2(new_n265_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n232_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT86), .B1(new_n266_), .B2(new_n232_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n271_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n268_), .A2(new_n270_), .A3(new_n232_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n276_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n280_), .B1(new_n283_), .B2(new_n271_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n275_), .A2(new_n280_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n278_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n279_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G1gat), .B(G29gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(G85gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT0), .B(G57gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n277_), .A2(KEYINPUT4), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n278_), .B1(new_n275_), .B2(new_n280_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n292_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n288_), .A2(new_n292_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298_));
  INV_X1    g097(.A(G197gat), .ZN(new_n299_));
  INV_X1    g098(.A(G204gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G197gat), .A2(G204gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(KEYINPUT21), .A3(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G211gat), .B(G218gat), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT21), .ZN(new_n306_));
  INV_X1    g105(.A(new_n302_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(G197gat), .A2(G204gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n204_), .A2(new_n207_), .B1(new_n213_), .B2(new_n211_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n205_), .A2(KEYINPUT25), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G183gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n206_), .A2(KEYINPUT26), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT26), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G190gat), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .A4(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(new_n223_), .A3(new_n224_), .A4(new_n204_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n312_), .B1(new_n320_), .B2(KEYINPUT84), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n223_), .A2(new_n224_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT84), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n204_), .A4(new_n319_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n311_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n305_), .A2(new_n310_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT20), .B1(new_n226_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT19), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n325_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n226_), .B2(new_n326_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n321_), .A2(new_n311_), .A3(new_n324_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n329_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G8gat), .B(G36gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT18), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n331_), .A2(new_n335_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n333_), .A2(new_n334_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n330_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n321_), .A2(new_n324_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n326_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n225_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n312_), .B1(new_n346_), .B2(new_n219_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n332_), .B1(new_n347_), .B2(new_n311_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n329_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n341_), .B1(new_n343_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n298_), .B1(new_n340_), .B2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n311_), .A2(new_n320_), .A3(new_n215_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n333_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n329_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n345_), .A2(new_n330_), .A3(new_n348_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n341_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n339_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(KEYINPUT27), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n297_), .A2(new_n351_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G228gat), .A2(G233gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT82), .Z(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n268_), .A2(KEYINPUT29), .A3(new_n270_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(new_n326_), .ZN(new_n365_));
  AOI211_X1 g164(.A(new_n362_), .B(new_n311_), .C1(new_n266_), .C2(KEYINPUT29), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n369_));
  XOR2_X1   g168(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G78gat), .B(G106gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT83), .ZN(new_n374_));
  XOR2_X1   g173(.A(G22gat), .B(G50gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n369_), .A2(new_n370_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n369_), .A2(new_n370_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n377_), .B(new_n378_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n372_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n376_), .B1(new_n372_), .B2(new_n379_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n240_), .B1(new_n360_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n339_), .A2(KEYINPUT32), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n386_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n384_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  OAI22_X1  g189(.A1(new_n297_), .A2(new_n390_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n295_), .A2(KEYINPUT33), .A3(new_n296_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT85), .B1(new_n340_), .B2(new_n350_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n343_), .A2(new_n349_), .A3(new_n341_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n358_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n292_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n277_), .B2(new_n286_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n285_), .A2(new_n278_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n400_), .B1(new_n284_), .B2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n393_), .A2(new_n398_), .A3(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n279_), .B(new_n399_), .C1(new_n284_), .C2(new_n287_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT33), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT87), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT87), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n408_), .A3(new_n405_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n403_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n392_), .B1(new_n410_), .B2(KEYINPUT88), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n398_), .A2(new_n402_), .ZN(new_n412_));
  AOI211_X1 g211(.A(KEYINPUT87), .B(KEYINPUT33), .C1(new_n295_), .C2(new_n296_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n408_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n412_), .B(new_n393_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT88), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n383_), .B1(new_n411_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n297_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n419_), .A2(new_n239_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n359_), .A2(new_n351_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n382_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n418_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G85gat), .ZN(new_n428_));
  INV_X1    g227(.A(G92gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G85gat), .A2(G92gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G99gat), .A2(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT6), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n439_));
  INV_X1    g238(.A(G99gat), .ZN(new_n440_));
  INV_X1    g239(.A(G106gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n433_), .B1(new_n438_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT8), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n436_), .B1(G99gat), .B2(G106gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n434_), .A2(KEYINPUT6), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n443_), .B(new_n442_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT8), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n433_), .ZN(new_n451_));
  OR2_X1    g250(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n441_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(KEYINPUT64), .A3(new_n441_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n435_), .A2(new_n437_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n430_), .A2(KEYINPUT9), .A3(new_n431_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n431_), .A2(KEYINPUT9), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n446_), .A2(new_n451_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G57gat), .B(G64gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G71gat), .B(G78gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(KEYINPUT11), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(KEYINPUT11), .ZN(new_n470_));
  INV_X1    g269(.A(new_n468_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n467_), .A2(KEYINPUT11), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n469_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n466_), .A2(KEYINPUT65), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n461_), .A2(new_n465_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n443_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI211_X1 g278(.A(KEYINPUT8), .B(new_n432_), .C1(new_n479_), .C2(new_n462_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n450_), .B1(new_n449_), .B2(new_n433_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n474_), .B(new_n476_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT65), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n476_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n474_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n475_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G230gat), .A2(G233gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT66), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT67), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n480_), .A2(new_n481_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT67), .B1(new_n446_), .B2(new_n451_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n476_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n486_), .A2(KEYINPUT12), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT12), .B1(new_n485_), .B2(new_n486_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n482_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n499_), .A2(new_n502_), .A3(new_n489_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT66), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n488_), .A2(new_n504_), .A3(new_n490_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n492_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G120gat), .B(G148gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT5), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G176gat), .B(G204gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n510_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n492_), .A2(new_n503_), .A3(new_n505_), .A4(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n511_), .A2(KEYINPUT13), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT13), .B1(new_n511_), .B2(new_n513_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G36gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(G29gat), .ZN(new_n519_));
  INV_X1    g318(.A(G29gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G36gat), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT68), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n521_), .A3(KEYINPUT68), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G43gat), .B(G50gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n525_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n519_), .A2(new_n521_), .A3(KEYINPUT68), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(new_n528_), .B2(new_n522_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G1gat), .B(G8gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(G22gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT72), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(G15gat), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n235_), .A2(KEYINPUT72), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n533_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n235_), .A2(KEYINPUT72), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(G15gat), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(G22gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT14), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(G1gat), .B2(G8gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n532_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  AOI211_X1 g344(.A(new_n531_), .B(new_n543_), .C1(new_n537_), .C2(new_n540_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n530_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n538_), .A2(new_n539_), .A3(G22gat), .ZN(new_n548_));
  AOI21_X1  g347(.A(G22gat), .B1(new_n538_), .B2(new_n539_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n544_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n531_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n532_), .B(new_n544_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n551_), .A2(new_n526_), .A3(new_n529_), .A4(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT74), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n551_), .A2(new_n552_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT74), .A3(new_n530_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n555_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT75), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT75), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n555_), .A2(new_n562_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT69), .B(KEYINPUT15), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n530_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n526_), .A2(new_n529_), .A3(new_n565_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n558_), .A3(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n569_), .A2(new_n556_), .A3(new_n553_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n564_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G113gat), .B(G141gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G169gat), .B(G197gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n564_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n517_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n427_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n558_), .B(new_n486_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G127gat), .B(G155gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT16), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT17), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n585_), .B1(new_n592_), .B2(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT73), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT73), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n591_), .A2(new_n596_), .A3(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT34), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT35), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(KEYINPUT35), .ZN(new_n602_));
  INV_X1    g401(.A(new_n530_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n466_), .B2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n601_), .B1(new_n604_), .B2(KEYINPUT70), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n493_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n446_), .A2(KEYINPUT67), .A3(new_n451_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n606_), .A2(new_n607_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n567_), .A2(new_n568_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n604_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n605_), .A2(new_n610_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G134gat), .B(G162gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT36), .Z(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n613_), .A2(KEYINPUT36), .A3(new_n617_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n617_), .A2(KEYINPUT36), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n614_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n618_), .B(KEYINPUT71), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n613_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n623_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n598_), .B1(new_n624_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n582_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT91), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT91), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n582_), .B2(new_n632_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n297_), .A2(G1gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT92), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n634_), .A2(KEYINPUT92), .A3(new_n636_), .A4(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n640_), .A2(KEYINPUT38), .A3(new_n641_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n413_), .A2(new_n414_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n416_), .B1(new_n646_), .B2(new_n403_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n403_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n648_), .B(KEYINPUT88), .C1(new_n414_), .C2(new_n413_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n649_), .A3(new_n392_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n425_), .B1(new_n650_), .B2(new_n383_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n622_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n598_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n516_), .A2(KEYINPUT93), .A3(new_n579_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT93), .B1(new_n516_), .B2(new_n579_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n652_), .A2(new_n653_), .A3(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n297_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT94), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n644_), .A2(new_n645_), .A3(new_n661_), .ZN(G1324gat));
  NOR2_X1   g461(.A1(new_n423_), .A2(G8gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n634_), .A2(new_n636_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n423_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n652_), .A2(new_n653_), .A3(new_n665_), .A4(new_n658_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT95), .B(KEYINPUT39), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(G8gat), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n666_), .B2(G8gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n664_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(KEYINPUT96), .B(KEYINPUT40), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n659_), .B2(new_n239_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT97), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT97), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(KEYINPUT41), .A3(new_n676_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n633_), .A2(new_n235_), .A3(new_n240_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(G1326gat));
  OAI21_X1  g481(.A(G22gat), .B1(new_n659_), .B2(new_n424_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT42), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n633_), .A2(new_n533_), .A3(new_n382_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(new_n622_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n653_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n383_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n391_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(new_n649_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n581_), .B(new_n688_), .C1(new_n691_), .C2(new_n425_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT99), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n427_), .A2(new_n694_), .A3(new_n581_), .A4(new_n688_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G29gat), .B1(new_n696_), .B2(new_n419_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n620_), .A2(new_n621_), .A3(KEYINPUT37), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(new_n629_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n700_), .B2(KEYINPUT98), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n624_), .A2(new_n630_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n651_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT98), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n700_), .B(new_n705_), .C1(new_n691_), .C2(new_n425_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n598_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT44), .B1(new_n707_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n711_), .B(new_n708_), .C1(new_n703_), .C2(new_n706_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n297_), .A2(new_n520_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n697_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(KEYINPUT46), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n423_), .A2(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n693_), .A2(new_n695_), .A3(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT100), .B(KEYINPUT45), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT101), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n721_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n693_), .A2(new_n695_), .A3(new_n723_), .A4(new_n718_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n717_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n716_), .A2(KEYINPUT46), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n710_), .A2(new_n712_), .A3(new_n423_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n725_), .B(new_n726_), .C1(new_n727_), .C2(new_n518_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n705_), .B1(new_n427_), .B2(new_n700_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n651_), .A2(new_n702_), .A3(new_n701_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n709_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n711_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n707_), .A2(KEYINPUT44), .A3(new_n709_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n665_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G36gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n726_), .B1(new_n736_), .B2(new_n725_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n729_), .A2(new_n737_), .ZN(G1329gat));
  NAND3_X1  g537(.A1(new_n713_), .A2(G43gat), .A3(new_n240_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n696_), .A2(new_n240_), .ZN(new_n740_));
  INV_X1    g539(.A(G43gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n739_), .A2(new_n742_), .A3(new_n744_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1330gat));
  INV_X1    g547(.A(G50gat), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n382_), .A2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT104), .Z(new_n751_));
  NAND2_X1  g550(.A1(new_n696_), .A2(new_n751_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n710_), .A2(new_n712_), .A3(new_n424_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n749_), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n516_), .A2(new_n579_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n653_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n652_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(G57gat), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n297_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(KEYINPUT105), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(KEYINPUT105), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n651_), .A2(new_n579_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n632_), .A2(new_n516_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G57gat), .B1(new_n766_), .B2(new_n419_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n762_), .A2(new_n763_), .A3(new_n767_), .ZN(G1332gat));
  NAND3_X1  g567(.A1(new_n652_), .A2(new_n665_), .A3(new_n757_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT48), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(G64gat), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n769_), .B2(G64gat), .ZN(new_n773_));
  INV_X1    g572(.A(new_n766_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n423_), .A2(G64gat), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT106), .ZN(new_n776_));
  OAI22_X1  g575(.A1(new_n772_), .A2(new_n773_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT107), .Z(G1333gat));
  NAND3_X1  g577(.A1(new_n652_), .A2(new_n240_), .A3(new_n757_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(G71gat), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n779_), .B2(G71gat), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n239_), .A2(G71gat), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT108), .Z(new_n785_));
  OAI22_X1  g584(.A1(new_n782_), .A2(new_n783_), .B1(new_n774_), .B2(new_n785_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT109), .Z(G1334gat));
  OAI21_X1  g586(.A(G78gat), .B1(new_n758_), .B2(new_n424_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT50), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n424_), .A2(G78gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n789_), .B1(new_n774_), .B2(new_n790_), .ZN(G1335gat));
  NAND3_X1  g590(.A1(new_n764_), .A2(new_n517_), .A3(new_n688_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n428_), .A3(new_n419_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n755_), .A2(new_n598_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n707_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT110), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n795_), .B1(new_n703_), .B2(new_n706_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n297_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n794_), .B1(new_n802_), .B2(new_n428_), .ZN(G1336gat));
  NAND3_X1  g602(.A1(new_n793_), .A2(new_n429_), .A3(new_n665_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n423_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n429_), .ZN(G1337gat));
  NAND3_X1  g605(.A1(new_n793_), .A2(new_n459_), .A3(new_n240_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n239_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n440_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(KEYINPUT111), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  OAI221_X1 g611(.A(new_n807_), .B1(KEYINPUT111), .B2(new_n810_), .C1(new_n808_), .C2(new_n440_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1338gat));
  NAND3_X1  g613(.A1(new_n793_), .A2(new_n441_), .A3(new_n382_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n799_), .A2(new_n382_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817_));
  OAI21_X1  g616(.A(G106gat), .B1(new_n817_), .B2(KEYINPUT112), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n816_), .A2(new_n819_), .B1(KEYINPUT112), .B2(new_n817_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(KEYINPUT112), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n821_), .B(new_n818_), .C1(new_n799_), .C2(new_n382_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n815_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT53), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n815_), .C1(new_n820_), .C2(new_n822_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1339gat));
  NAND2_X1  g626(.A1(new_n424_), .A2(new_n423_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n828_), .A2(new_n297_), .A3(new_n239_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT12), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n466_), .B2(new_n474_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n482_), .C1(new_n608_), .C2(new_n497_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n835_), .B2(new_n490_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n490_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n499_), .A2(new_n502_), .A3(KEYINPUT55), .A4(new_n489_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n831_), .B(new_n510_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n513_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n489_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n503_), .B1(new_n843_), .B2(new_n832_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n839_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n831_), .B1(new_n845_), .B2(new_n510_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n842_), .A2(new_n580_), .A3(new_n846_), .ZN(new_n847_));
  AOI211_X1 g646(.A(new_n570_), .B(new_n576_), .C1(new_n561_), .C2(new_n563_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n553_), .A2(new_n557_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n575_), .B1(new_n849_), .B2(new_n569_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n555_), .A2(new_n556_), .A3(new_n559_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT113), .B1(new_n848_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n578_), .A2(new_n855_), .A3(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n511_), .A2(new_n513_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n687_), .B1(new_n847_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n513_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n512_), .B1(new_n844_), .B2(new_n839_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n831_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n510_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT56), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n579_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n859_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(KEYINPUT57), .A3(new_n687_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n863_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n866_), .A2(new_n868_), .A3(new_n857_), .A4(KEYINPUT114), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT115), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n866_), .A2(new_n857_), .A3(new_n868_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT114), .B1(new_n878_), .B2(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n702_), .B1(new_n876_), .B2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n598_), .B1(new_n872_), .B2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n653_), .B(new_n580_), .C1(new_n629_), .C2(new_n699_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n883_), .B2(new_n517_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n631_), .A2(new_n885_), .A3(new_n516_), .A4(new_n580_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n830_), .B1(new_n882_), .B2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G113gat), .B1(new_n888_), .B2(new_n579_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n870_), .B2(new_n687_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n862_), .B(new_n622_), .C1(new_n869_), .C2(new_n859_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n880_), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT58), .B1(new_n873_), .B2(KEYINPUT115), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n700_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n653_), .B1(new_n894_), .B2(new_n897_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n884_), .A2(new_n886_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n891_), .B1(new_n900_), .B2(new_n830_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n829_), .B(new_n903_), .C1(new_n898_), .C2(new_n899_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n901_), .A2(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT117), .B(G113gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n579_), .A2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT118), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n889_), .B1(new_n905_), .B2(new_n908_), .ZN(G1340gat));
  OAI211_X1 g708(.A(new_n517_), .B(new_n904_), .C1(new_n888_), .C2(new_n890_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT119), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n516_), .B2(G120gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n888_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n901_), .A2(new_n915_), .A3(new_n517_), .A4(new_n904_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n911_), .A2(new_n914_), .A3(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G120gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n888_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1341gat));
  INV_X1    g719(.A(G127gat), .ZN(new_n921_));
  INV_X1    g720(.A(new_n888_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n598_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n923_), .A2(KEYINPUT120), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n905_), .A2(G127gat), .A3(new_n653_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(KEYINPUT120), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .ZN(G1342gat));
  NAND2_X1  g726(.A1(new_n905_), .A2(new_n700_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(G134gat), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n687_), .A2(G134gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n922_), .B2(new_n930_), .ZN(G1343gat));
  NAND2_X1  g730(.A1(new_n882_), .A2(new_n887_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n424_), .A2(new_n240_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n665_), .A2(new_n297_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n580_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(new_n248_), .ZN(G1344gat));
  NOR2_X1   g736(.A1(new_n935_), .A2(new_n516_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n249_), .ZN(G1345gat));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n940_), .B1(new_n935_), .B2(new_n598_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n933_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n900_), .A2(new_n942_), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n943_), .A2(KEYINPUT121), .A3(new_n653_), .A4(new_n934_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n941_), .A2(new_n944_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(KEYINPUT61), .B(G155gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(G1346gat));
  OAI21_X1  g746(.A(G162gat), .B1(new_n935_), .B2(new_n702_), .ZN(new_n948_));
  OR2_X1    g747(.A1(new_n687_), .A2(G162gat), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n935_), .B2(new_n949_), .ZN(G1347gat));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n665_), .A2(new_n424_), .A3(new_n420_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n900_), .B2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n952_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n932_), .A2(KEYINPUT122), .A3(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n953_), .A2(new_n955_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(KEYINPUT22), .B(G169gat), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n956_), .A2(new_n579_), .A3(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n900_), .A2(new_n952_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n579_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n959_), .B1(new_n961_), .B2(G169gat), .ZN(new_n962_));
  AOI211_X1 g761(.A(KEYINPUT62), .B(new_n212_), .C1(new_n960_), .C2(new_n579_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n958_), .B1(new_n962_), .B2(new_n963_), .ZN(G1348gat));
  NAND2_X1  g763(.A1(new_n517_), .A2(new_n210_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n965_), .B1(new_n953_), .B2(new_n955_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n210_), .B1(new_n960_), .B2(new_n517_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n968_));
  OR3_X1    g767(.A1(new_n966_), .A2(new_n967_), .A3(new_n968_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n968_), .B1(new_n966_), .B2(new_n967_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1349gat));
  AOI21_X1  g770(.A(G183gat), .B1(new_n960_), .B2(new_n653_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n598_), .A2(new_n217_), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n972_), .B1(new_n956_), .B2(new_n973_), .ZN(G1350gat));
  INV_X1    g773(.A(new_n956_), .ZN(new_n975_));
  OAI21_X1  g774(.A(G190gat), .B1(new_n975_), .B2(new_n702_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n622_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n975_), .B2(new_n977_), .ZN(G1351gat));
  NOR2_X1   g777(.A1(new_n423_), .A2(new_n419_), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n932_), .A2(new_n933_), .A3(new_n979_), .ZN(new_n980_));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n980_), .A2(new_n981_), .ZN(new_n982_));
  NAND4_X1  g781(.A1(new_n932_), .A2(KEYINPUT124), .A3(new_n933_), .A4(new_n979_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n982_), .A2(new_n983_), .ZN(new_n984_));
  OR2_X1    g783(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n985_));
  AND3_X1   g784(.A1(new_n984_), .A2(new_n579_), .A3(new_n985_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n987_));
  AOI22_X1  g786(.A1(new_n984_), .A2(new_n579_), .B1(new_n987_), .B2(new_n985_), .ZN(new_n988_));
  NOR2_X1   g787(.A1(new_n986_), .A2(new_n988_), .ZN(G1352gat));
  AOI21_X1  g788(.A(new_n516_), .B1(new_n982_), .B2(new_n983_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(new_n990_), .B(new_n300_), .ZN(G1353gat));
  AOI21_X1  g790(.A(new_n598_), .B1(new_n982_), .B2(new_n983_), .ZN(new_n992_));
  NOR2_X1   g791(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n993_));
  AND2_X1   g792(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n992_), .B1(new_n993_), .B2(new_n994_), .ZN(new_n995_));
  OAI21_X1  g794(.A(new_n995_), .B1(new_n992_), .B2(new_n993_), .ZN(G1354gat));
  NAND2_X1  g795(.A1(new_n984_), .A2(new_n622_), .ZN(new_n997_));
  XOR2_X1   g796(.A(KEYINPUT126), .B(G218gat), .Z(new_n998_));
  NOR2_X1   g797(.A1(new_n702_), .A2(new_n998_), .ZN(new_n999_));
  AOI22_X1  g798(.A1(new_n997_), .A2(new_n998_), .B1(new_n984_), .B2(new_n999_), .ZN(G1355gat));
endmodule


