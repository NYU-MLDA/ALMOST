//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  AND2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(G141gat), .ZN(new_n205_));
  INV_X1    g004(.A(G148gat), .ZN(new_n206_));
  AOI22_X1  g005(.A1(new_n204_), .A2(KEYINPUT1), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G155gat), .B(G162gat), .ZN(new_n208_));
  OAI221_X1 g007(.A(new_n207_), .B1(new_n205_), .B2(new_n206_), .C1(KEYINPUT1), .C2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(KEYINPUT90), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NOR3_X1   g011(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n215_));
  NOR4_X1   g014(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n209_), .B1(new_n210_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT29), .ZN(new_n218_));
  INV_X1    g017(.A(G228gat), .ZN(new_n219_));
  INV_X1    g018(.A(G233gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT21), .ZN(new_n224_));
  OR3_X1    g023(.A1(new_n223_), .A2(KEYINPUT92), .A3(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G211gat), .B(G218gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n224_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT92), .B1(new_n223_), .B2(new_n224_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n226_), .A2(KEYINPUT93), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n223_), .A2(new_n224_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(KEYINPUT93), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n218_), .A2(new_n222_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n222_), .B1(new_n218_), .B2(new_n234_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n203_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT95), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n237_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(new_n235_), .A3(new_n202_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT94), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT94), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n241_), .A2(new_n244_), .A3(new_n235_), .A4(new_n202_), .ZN(new_n245_));
  OAI211_X1 g044(.A(KEYINPUT95), .B(new_n203_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n240_), .A2(new_n243_), .A3(new_n245_), .A4(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n217_), .A2(KEYINPUT29), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G22gat), .B(G50gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n248_), .B(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT96), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n242_), .B2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n255_), .B(new_n238_), .C1(new_n254_), .C2(new_n242_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT89), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT30), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT22), .B(G169gat), .ZN(new_n260_));
  INV_X1    g059(.A(G176gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT88), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT23), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT87), .B(G183gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(new_n269_), .B2(G190gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT88), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n262_), .A2(new_n271_), .A3(new_n263_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G190gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT25), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n268_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n274_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G169gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n261_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n280_), .A2(KEYINPUT24), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(KEYINPUT24), .A3(new_n263_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n278_), .A2(new_n281_), .A3(new_n282_), .A4(new_n267_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n259_), .B1(new_n273_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G113gat), .B(G120gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(G127gat), .B(G134gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n273_), .A2(new_n283_), .A3(new_n259_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n285_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n290_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n288_), .B1(new_n292_), .B2(new_n284_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G43gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT31), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n296_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G71gat), .B(G99gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G227gat), .A2(G233gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n298_), .A2(new_n299_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n291_), .A2(new_n293_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n295_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n306_), .B2(new_n297_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n258_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n303_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n302_), .A3(new_n297_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT89), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n257_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n310_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n253_), .A3(new_n256_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n217_), .B(new_n289_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT4), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT4), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n217_), .A2(new_n320_), .A3(new_n288_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(new_n318_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G1gat), .B(G29gat), .ZN(new_n325_));
  INV_X1    g124(.A(G85gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT0), .B(G57gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n322_), .A2(new_n323_), .A3(new_n329_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n273_), .A2(new_n283_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n234_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n267_), .B1(G183gat), .B2(G190gat), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n263_), .A2(KEYINPUT98), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n263_), .A2(KEYINPUT98), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n336_), .A2(new_n262_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n280_), .A2(new_n263_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT25), .B(G183gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n274_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n279_), .A3(new_n261_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n342_), .A2(new_n267_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n339_), .A2(new_n229_), .A3(new_n233_), .A4(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n335_), .A2(KEYINPUT20), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT19), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n339_), .A2(new_n346_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n234_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(KEYINPUT20), .C1(new_n234_), .C2(new_n334_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n351_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G8gat), .B(G36gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n360_), .B(KEYINPUT104), .Z(new_n361_));
  NAND3_X1  g160(.A1(new_n355_), .A2(KEYINPUT105), .A3(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n347_), .A2(KEYINPUT99), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT20), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n347_), .B2(KEYINPUT99), .ZN(new_n365_));
  INV_X1    g164(.A(new_n350_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n363_), .A2(new_n365_), .A3(new_n366_), .A4(new_n335_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n354_), .A2(new_n350_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n360_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n362_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT105), .B1(new_n355_), .B2(new_n361_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT27), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT101), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n367_), .A2(new_n368_), .A3(KEYINPUT101), .A4(new_n369_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n367_), .A2(new_n368_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT102), .B1(new_n379_), .B2(new_n360_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n379_), .A2(KEYINPUT102), .A3(new_n360_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n377_), .B(new_n378_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n333_), .B1(new_n373_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n315_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n369_), .A2(KEYINPUT32), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n355_), .A2(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n333_), .B(new_n387_), .C1(new_n379_), .C2(new_n386_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n316_), .A2(new_n319_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n330_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n390_), .A2(KEYINPUT103), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n317_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(KEYINPUT103), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n377_), .B(new_n394_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n332_), .B(KEYINPUT33), .Z(new_n396_));
  OAI21_X1  g195(.A(new_n388_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n257_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n308_), .A2(new_n311_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n384_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G230gat), .A2(G233gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n402_), .B(KEYINPUT64), .Z(new_n403_));
  INV_X1    g202(.A(KEYINPUT69), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n326_), .A2(G92gat), .ZN(new_n405_));
  INV_X1    g204(.A(G92gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(G85gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(G85gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n326_), .A2(G92gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(KEYINPUT69), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G99gat), .A2(G106gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT71), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT6), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(KEYINPUT71), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n414_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(KEYINPUT71), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(KEYINPUT6), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n413_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n419_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NOR4_X1   g223(.A1(KEYINPUT68), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT68), .ZN(new_n426_));
  NOR2_X1   g225(.A1(G99gat), .A2(G106gat), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT7), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n412_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT8), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n417_), .A2(G99gat), .A3(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n435_), .B(new_n423_), .C1(new_n425_), .C2(new_n429_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT8), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n412_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT70), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n436_), .A2(new_n412_), .A3(KEYINPUT70), .A4(new_n437_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n432_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(KEYINPUT10), .B(G99gat), .Z(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT65), .B(G106gat), .Z(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT66), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n446_), .A2(new_n326_), .A3(KEYINPUT9), .ZN(new_n447_));
  NOR2_X1   g246(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(G92gat), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT9), .B1(new_n405_), .B2(new_n407_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n445_), .A2(new_n449_), .A3(new_n450_), .A4(new_n435_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT67), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n442_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G57gat), .B(G64gat), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n454_), .A2(KEYINPUT11), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(KEYINPUT11), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G71gat), .B(G78gat), .ZN(new_n457_));
  OR3_X1    g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n457_), .A3(KEYINPUT11), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n453_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n442_), .A2(new_n452_), .A3(new_n460_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(KEYINPUT12), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n460_), .B1(new_n442_), .B2(new_n452_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT12), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n403_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n403_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G120gat), .B(G148gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(G204gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT5), .B(G176gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(KEYINPUT72), .ZN(new_n476_));
  OR3_X1    g275(.A1(new_n468_), .A2(new_n470_), .A3(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT13), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(KEYINPUT13), .A3(new_n478_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT81), .B(G1gat), .Z(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G1gat), .B(G8gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT74), .B(G43gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G29gat), .ZN(new_n492_));
  INV_X1    g291(.A(G36gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G50gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G29gat), .A2(G36gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n491_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(new_n490_), .A3(new_n497_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n489_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n500_), .A2(new_n502_), .A3(KEYINPUT15), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  MUX2_X1   g311(.A(new_n504_), .B(new_n512_), .S(new_n489_), .Z(new_n513_));
  AOI21_X1  g312(.A(new_n508_), .B1(new_n506_), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515_));
  INV_X1    g314(.A(G197gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT86), .B(G169gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT85), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n514_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n482_), .A2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n401_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G231gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n460_), .B(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n527_), .B(new_n489_), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT84), .B(G127gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G183gat), .B(G211gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G155gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n532_), .B(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(KEYINPUT82), .A3(KEYINPUT17), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(KEYINPUT17), .B2(new_n535_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n529_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n528_), .A2(new_n536_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT79), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n442_), .A2(new_n503_), .A3(new_n452_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n512_), .B1(new_n442_), .B2(new_n452_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT75), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT75), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n453_), .B2(new_n504_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT35), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n544_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT78), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n544_), .A2(new_n546_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n544_), .A2(KEYINPUT78), .A3(new_n546_), .A4(new_n550_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n553_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  INV_X1    g359(.A(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT76), .B(G190gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT36), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT77), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n553_), .A2(new_n557_), .A3(new_n558_), .A4(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n541_), .B1(new_n566_), .B2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n541_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT37), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT80), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n566_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n559_), .A2(KEYINPUT80), .A3(new_n565_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n570_), .A4(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n525_), .A2(new_n540_), .A3(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n333_), .A3(new_n483_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT38), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n575_), .A2(new_n570_), .A3(new_n577_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n401_), .A2(KEYINPUT107), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT107), .B1(new_n401_), .B2(new_n583_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n540_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n524_), .A2(KEYINPUT106), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n524_), .A2(KEYINPUT106), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n333_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n582_), .A2(new_n593_), .ZN(G1324gat));
  NAND2_X1  g393(.A1(new_n373_), .A2(new_n382_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n587_), .A2(new_n590_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(G8gat), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(KEYINPUT108), .A3(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n580_), .A2(new_n484_), .A3(new_n596_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n599_), .A2(KEYINPUT108), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(KEYINPUT108), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n597_), .A2(G8gat), .A3(new_n602_), .A4(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n600_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g405(.A(G15gat), .B1(new_n591_), .B2(new_n399_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT41), .Z(new_n608_));
  INV_X1    g407(.A(G15gat), .ZN(new_n609_));
  INV_X1    g408(.A(new_n399_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n580_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(G1326gat));
  OAI21_X1  g411(.A(G22gat), .B1(new_n591_), .B2(new_n398_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT42), .ZN(new_n614_));
  INV_X1    g413(.A(G22gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n580_), .A2(new_n615_), .A3(new_n257_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(G1327gat));
  NOR2_X1   g416(.A1(new_n583_), .A2(new_n540_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n525_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(G29gat), .B1(new_n620_), .B2(new_n333_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n401_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT43), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT109), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n623_), .A2(KEYINPUT43), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT109), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n627_), .A3(KEYINPUT43), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n626_), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n540_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n622_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n631_), .A2(new_n492_), .A3(new_n592_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(KEYINPUT44), .A3(new_n630_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n621_), .B1(new_n632_), .B2(new_n633_), .ZN(G1328gat));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n596_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT111), .B1(new_n635_), .B2(new_n631_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n631_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT111), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n596_), .A4(new_n633_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n636_), .A2(new_n639_), .A3(G36gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n620_), .A2(new_n493_), .A3(new_n596_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT45), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT46), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(KEYINPUT46), .A3(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1329gat));
  NAND3_X1  g446(.A1(new_n633_), .A2(G43gat), .A3(new_n313_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n619_), .A2(new_n399_), .ZN(new_n649_));
  OAI22_X1  g448(.A1(new_n648_), .A2(new_n631_), .B1(G43gat), .B2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(G1330gat));
  NAND3_X1  g451(.A1(new_n620_), .A2(new_n495_), .A3(new_n257_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n637_), .A2(new_n257_), .A3(new_n633_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT113), .A3(G50gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT113), .B1(new_n654_), .B2(G50gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(G1331gat));
  INV_X1    g456(.A(new_n482_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n522_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n587_), .A2(G57gat), .A3(new_n333_), .A4(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT115), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n579_), .A2(new_n482_), .A3(new_n540_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT114), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n522_), .B1(new_n384_), .B2(new_n400_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(KEYINPUT114), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G57gat), .B1(new_n666_), .B2(new_n333_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n661_), .A2(new_n667_), .ZN(G1332gat));
  NAND2_X1  g467(.A1(new_n587_), .A2(new_n659_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G64gat), .B1(new_n669_), .B2(new_n595_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT48), .ZN(new_n671_));
  INV_X1    g470(.A(G64gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n672_), .A3(new_n596_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(G1333gat));
  OAI21_X1  g473(.A(G71gat), .B1(new_n669_), .B2(new_n399_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT49), .ZN(new_n676_));
  INV_X1    g475(.A(G71gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n666_), .A2(new_n677_), .A3(new_n610_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1334gat));
  OAI21_X1  g478(.A(G78gat), .B1(new_n669_), .B2(new_n398_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT50), .ZN(new_n681_));
  INV_X1    g480(.A(G78gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n666_), .A2(new_n682_), .A3(new_n257_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1335gat));
  NAND3_X1  g483(.A1(new_n664_), .A2(new_n618_), .A3(new_n482_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G85gat), .B1(new_n686_), .B2(new_n333_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n629_), .A2(new_n586_), .A3(new_n659_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n446_), .A2(new_n326_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n333_), .B1(new_n448_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT116), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n687_), .B1(new_n688_), .B2(new_n691_), .ZN(G1336gat));
  AOI21_X1  g491(.A(G92gat), .B1(new_n686_), .B2(new_n596_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n595_), .A2(new_n406_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n688_), .B2(new_n694_), .ZN(G1337gat));
  NAND3_X1  g494(.A1(new_n686_), .A2(new_n443_), .A3(new_n313_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n688_), .A2(new_n610_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT117), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(G99gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n697_), .B2(G99gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT51), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(KEYINPUT118), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  OAI221_X1 g503(.A(new_n696_), .B1(KEYINPUT118), .B2(new_n702_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1338gat));
  NAND3_X1  g505(.A1(new_n686_), .A2(new_n444_), .A3(new_n257_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n688_), .A2(new_n257_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT52), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G106gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G106gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT53), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT53), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n707_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1339gat));
  INV_X1    g515(.A(new_n314_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n596_), .A2(new_n592_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n482_), .A2(new_n522_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n579_), .A2(new_n540_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT119), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT119), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n579_), .A2(new_n722_), .A3(new_n540_), .A4(new_n719_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n721_), .A2(KEYINPUT54), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT54), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n720_), .A2(KEYINPUT119), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n464_), .A2(new_n403_), .A3(new_n467_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n442_), .A2(new_n460_), .A3(new_n452_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n730_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n467_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n469_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT55), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n468_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n729_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT56), .B1(new_n737_), .B2(new_n475_), .ZN(new_n738_));
  MUX2_X1   g537(.A(new_n505_), .B(new_n513_), .S(new_n507_), .Z(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(new_n520_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n520_), .B2(new_n514_), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n468_), .A2(new_n470_), .A3(new_n474_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n464_), .A2(new_n467_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n735_), .B1(new_n743_), .B2(new_n469_), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT55), .B(new_n403_), .C1(new_n464_), .C2(new_n467_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n728_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n474_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n738_), .A2(new_n741_), .A3(new_n742_), .A4(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT121), .B1(new_n751_), .B2(new_n579_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT58), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n749_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n749_), .A2(new_n750_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT121), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n573_), .A4(new_n578_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n752_), .A2(new_n754_), .A3(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n738_), .A2(new_n522_), .A3(new_n742_), .A4(new_n748_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n477_), .A2(new_n478_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n741_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n762_), .A2(KEYINPUT57), .A3(new_n583_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT57), .B1(new_n762_), .B2(new_n583_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n540_), .B1(new_n758_), .B2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n717_), .B(new_n718_), .C1(new_n727_), .C2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G113gat), .B1(new_n768_), .B2(new_n522_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n724_), .A2(new_n726_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n758_), .A2(new_n765_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n586_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n773_), .A2(new_n717_), .A3(new_n718_), .A4(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT122), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(KEYINPUT59), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n767_), .A2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n775_), .A2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n779_), .A2(new_n523_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n769_), .B1(new_n780_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g580(.A(G120gat), .B1(new_n779_), .B2(new_n658_), .ZN(new_n782_));
  INV_X1    g581(.A(G120gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n658_), .B2(KEYINPUT60), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT60), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(KEYINPUT123), .B2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n768_), .B(new_n786_), .C1(KEYINPUT123), .C2(new_n784_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n782_), .A2(new_n787_), .ZN(G1341gat));
  AOI21_X1  g587(.A(G127gat), .B1(new_n768_), .B2(new_n540_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n779_), .A2(new_n586_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g590(.A(G134gat), .ZN(new_n792_));
  INV_X1    g591(.A(new_n583_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n768_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n579_), .B1(new_n775_), .B2(new_n778_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT124), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT124), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n798_), .B(new_n794_), .C1(new_n795_), .C2(new_n792_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1343gat));
  AOI21_X1  g599(.A(new_n312_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n718_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n523_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(new_n205_), .ZN(G1344gat));
  NOR2_X1   g603(.A1(new_n802_), .A2(new_n658_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(new_n206_), .ZN(G1345gat));
  INV_X1    g605(.A(new_n802_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n540_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT61), .B(G155gat), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  INV_X1    g609(.A(G162gat), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n802_), .A2(new_n811_), .A3(new_n579_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n807_), .A2(new_n793_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(new_n813_), .ZN(G1347gat));
  NOR3_X1   g613(.A1(new_n399_), .A2(new_n595_), .A3(new_n333_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n773_), .A2(new_n398_), .A3(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G169gat), .B1(new_n816_), .B2(new_n523_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT125), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT125), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n819_), .B(G169gat), .C1(new_n816_), .C2(new_n523_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(KEYINPUT62), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n816_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n522_), .A3(new_n260_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT62), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n817_), .A2(KEYINPUT125), .A3(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(new_n823_), .A3(new_n825_), .ZN(G1348gat));
  OAI21_X1  g625(.A(new_n261_), .B1(new_n816_), .B2(new_n658_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n398_), .B1(new_n727_), .B2(new_n766_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT126), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT126), .B(new_n398_), .C1(new_n727_), .C2(new_n766_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n658_), .A2(new_n261_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n830_), .A2(new_n815_), .A3(new_n831_), .A4(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n827_), .A2(new_n833_), .ZN(G1349gat));
  NAND4_X1  g633(.A1(new_n830_), .A2(new_n540_), .A3(new_n815_), .A4(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n268_), .ZN(new_n836_));
  OR3_X1    g635(.A1(new_n816_), .A2(new_n586_), .A3(new_n343_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT127), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT127), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n836_), .A2(new_n837_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1350gat));
  OAI21_X1  g641(.A(G190gat), .B1(new_n816_), .B2(new_n579_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n793_), .A2(new_n274_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n816_), .B2(new_n844_), .ZN(G1351gat));
  NOR2_X1   g644(.A1(new_n595_), .A2(new_n333_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n801_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n523_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(new_n516_), .ZN(G1352gat));
  INV_X1    g648(.A(new_n847_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n482_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g651(.A(KEYINPUT63), .B(G211gat), .C1(new_n850_), .C2(new_n540_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT63), .B(G211gat), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n847_), .A2(new_n586_), .A3(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1354gat));
  NOR3_X1   g655(.A1(new_n847_), .A2(new_n561_), .A3(new_n579_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n850_), .A2(new_n793_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n561_), .B2(new_n858_), .ZN(G1355gat));
endmodule


