//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G155gat), .ZN(new_n203_));
  INV_X1    g002(.A(G162gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(KEYINPUT1), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  AND2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT86), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT86), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n208_), .B(new_n209_), .C1(new_n210_), .C2(KEYINPUT1), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n207_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G141gat), .ZN(new_n215_));
  INV_X1    g014(.A(G148gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT87), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(new_n206_), .B2(new_n210_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n203_), .A2(new_n204_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(KEYINPUT87), .A3(new_n209_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT2), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n226_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n221_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G127gat), .B(G134gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n238_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT4), .A3(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n240_), .A2(KEYINPUT4), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n239_), .A2(new_n240_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G1gat), .B(G29gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G85gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT0), .B(G57gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n249_), .B(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT74), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(KEYINPUT13), .ZN(new_n256_));
  XOR2_X1   g055(.A(G71gat), .B(G78gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(G57gat), .B(G64gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n257_), .B1(KEYINPUT11), .B2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT69), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n258_), .A2(KEYINPUT11), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  OR3_X1    g061(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G99gat), .A2(G106gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT6), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT8), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G85gat), .A2(G92gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G85gat), .A2(G92gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n268_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n263_), .B(new_n264_), .C1(new_n276_), .C2(new_n266_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT66), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT6), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n266_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n275_), .B(new_n273_), .C1(new_n277_), .C2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT8), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n283_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n276_), .A2(new_n266_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n265_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n275_), .B1(new_n289_), .B2(new_n273_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n274_), .B1(new_n286_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT10), .B(G99gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT64), .ZN(new_n294_));
  INV_X1    g093(.A(G106gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT9), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n270_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT65), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n272_), .B1(new_n271_), .B2(KEYINPUT9), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n296_), .A2(new_n301_), .A3(new_n267_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n291_), .A2(new_n292_), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n292_), .B1(new_n291_), .B2(new_n302_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n262_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT70), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n291_), .A2(new_n302_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT68), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n291_), .A2(new_n292_), .A3(new_n302_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(new_n262_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n262_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n308_), .A2(new_n309_), .A3(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n306_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G230gat), .ZN(new_n316_));
  INV_X1    g115(.A(G233gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n302_), .B(KEYINPUT71), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n291_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT12), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n262_), .A2(new_n324_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n314_), .A2(new_n321_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n318_), .B1(new_n310_), .B2(new_n262_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n319_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G120gat), .B(G148gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G176gat), .B(G204gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n319_), .A2(new_n328_), .A3(new_n334_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n256_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(new_n337_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n339_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n341_), .A2(new_n342_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT75), .B1(new_n345_), .B2(new_n338_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G29gat), .B(G36gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G43gat), .B(G50gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT15), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G15gat), .B(G22gat), .ZN(new_n352_));
  INV_X1    g151(.A(G8gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G1gat), .B(G8gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n350_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G229gat), .A2(G233gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n357_), .B(new_n359_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n361_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G113gat), .B(G141gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G169gat), .B(G197gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  OR2_X1    g168(.A1(new_n369_), .A2(KEYINPUT78), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n366_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G231gat), .A2(G233gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n357_), .B(new_n372_), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n262_), .B(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G127gat), .B(G155gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT16), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G183gat), .B(G211gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT17), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n378_), .A2(new_n379_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n374_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n374_), .A2(new_n380_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT35), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G232gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT34), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n323_), .A2(new_n351_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n310_), .A2(new_n350_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n390_), .A2(new_n387_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n391_), .B(new_n392_), .C1(new_n387_), .C2(new_n390_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT76), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G190gat), .B(G218gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(G134gat), .B(G162gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT36), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n401_), .A2(KEYINPUT36), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n397_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n404_), .ZN(new_n406_));
  AOI221_X4 g205(.A(KEYINPUT76), .B1(new_n406_), .B2(new_n402_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n386_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n397_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n395_), .A2(new_n396_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n402_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n409_), .A2(new_n412_), .A3(new_n406_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n407_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n408_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR4_X1   g217(.A1(new_n347_), .A2(new_n371_), .A3(new_n385_), .A4(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT101), .ZN(new_n420_));
  INV_X1    g219(.A(new_n254_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n214_), .A2(new_n220_), .B1(new_n226_), .B2(new_n233_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n209_), .B1(new_n210_), .B2(KEYINPUT1), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n212_), .B1(new_n426_), .B2(KEYINPUT86), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n219_), .B1(new_n427_), .B2(new_n211_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n233_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT88), .B(KEYINPUT29), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT21), .ZN(new_n431_));
  AND2_X1   g230(.A1(G197gat), .A2(G204gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G197gat), .A2(G204gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G197gat), .ZN(new_n435_));
  INV_X1    g234(.A(G204gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G197gat), .A2(G204gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(KEYINPUT21), .A3(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G211gat), .B(G218gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n434_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G218gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G211gat), .ZN(new_n443_));
  INV_X1    g242(.A(G211gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G218gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(KEYINPUT21), .A3(new_n437_), .A4(new_n438_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n441_), .A2(KEYINPUT90), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT90), .B1(new_n441_), .B2(new_n447_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G228gat), .A2(G233gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n450_), .B(KEYINPUT89), .Z(new_n451_));
  NOR3_X1   g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n425_), .A2(new_n430_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n441_), .A2(new_n447_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n451_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G22gat), .B(G50gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT28), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n461_));
  NOR4_X1   g260(.A1(new_n428_), .A2(new_n429_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n459_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n221_), .A2(new_n424_), .A3(new_n234_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT28), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n423_), .A2(new_n460_), .A3(new_n424_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n458_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n457_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n453_), .A2(new_n456_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(new_n467_), .A3(new_n463_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT92), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n470_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n473_), .B1(new_n457_), .B2(new_n468_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT93), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n469_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G78gat), .B(G106gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT91), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n477_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n477_), .B2(new_n481_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n421_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT22), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G169gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT80), .ZN(new_n489_));
  AOI21_X1  g288(.A(G176gat), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT22), .B(G169gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n490_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT81), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G183gat), .A2(G190gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(G183gat), .A2(G190gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT82), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n496_), .A2(new_n497_), .A3(KEYINPUT82), .A4(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G169gat), .A2(G176gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT81), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n490_), .B(new_n505_), .C1(new_n489_), .C2(new_n491_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n493_), .A2(new_n503_), .A3(new_n504_), .A4(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n496_), .A2(new_n498_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n509_));
  NOR2_X1   g308(.A1(G169gat), .A2(G176gat), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT26), .B(G190gat), .ZN(new_n512_));
  INV_X1    g311(.A(G183gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT25), .B1(new_n513_), .B2(KEYINPUT79), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(KEYINPUT25), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n512_), .B(new_n514_), .C1(new_n515_), .C2(KEYINPUT79), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n504_), .A2(KEYINPUT24), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n511_), .B(new_n516_), .C1(new_n510_), .C2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT83), .B1(new_n507_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n507_), .A2(KEYINPUT83), .A3(new_n518_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n448_), .A2(new_n449_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT20), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n510_), .B1(new_n517_), .B2(KEYINPUT96), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(KEYINPUT96), .B2(new_n517_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT25), .B(G183gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n512_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n511_), .A3(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n504_), .B(KEYINPUT97), .Z(new_n531_));
  INV_X1    g330(.A(G176gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n491_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n499_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n525_), .B1(new_n535_), .B2(new_n454_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n524_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G226gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT95), .ZN(new_n539_));
  XOR2_X1   g338(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G8gat), .B(G36gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G64gat), .B(G92gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n521_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n522_), .B1(new_n549_), .B2(new_n519_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n530_), .A2(new_n441_), .A3(new_n447_), .A4(new_n534_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n551_), .A2(KEYINPUT20), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n541_), .A3(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n543_), .A2(new_n548_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n548_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n541_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n520_), .A2(new_n521_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n522_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n541_), .B1(new_n524_), .B2(new_n536_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n555_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n560_), .A3(KEYINPUT99), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT27), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT99), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n563_), .B(new_n555_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n537_), .A2(new_n542_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n552_), .B(KEYINPUT100), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n550_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n566_), .B1(new_n568_), .B2(new_n542_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT27), .B(new_n554_), .C1(new_n569_), .C2(new_n548_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n420_), .B1(new_n486_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n477_), .A2(new_n481_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n483_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n477_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n565_), .A2(new_n570_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT101), .A4(new_n421_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n561_), .A2(new_n564_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n249_), .A2(new_n253_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT33), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n249_), .A2(KEYINPUT33), .A3(new_n253_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n247_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n253_), .B1(new_n585_), .B2(new_n245_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n245_), .B2(new_n243_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n580_), .A2(new_n583_), .A3(new_n584_), .A4(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n548_), .A2(KEYINPUT32), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n543_), .A2(new_n553_), .A3(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n254_), .B(new_n590_), .C1(new_n569_), .C2(new_n589_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n484_), .A2(new_n485_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n572_), .A2(new_n579_), .A3(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G15gat), .B(G43gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(G71gat), .B(G99gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n557_), .B(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G227gat), .A2(G233gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT84), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT30), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n602_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT85), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(KEYINPUT85), .A3(new_n604_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n605_), .A2(new_n606_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n595_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT102), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n613_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n577_), .A2(new_n571_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n421_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n595_), .A2(KEYINPUT102), .A3(new_n613_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n419_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT103), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n419_), .A2(new_n624_), .A3(new_n621_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n623_), .A2(KEYINPUT104), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT104), .B1(new_n623_), .B2(new_n625_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n202_), .B(new_n254_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n405_), .A2(new_n407_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n621_), .A2(KEYINPUT105), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT105), .B1(new_n621_), .B2(new_n631_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n347_), .A2(new_n371_), .A3(new_n385_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n254_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G1gat), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n628_), .A2(new_n629_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n630_), .A2(new_n637_), .A3(new_n638_), .ZN(G1324gat));
  OAI211_X1 g438(.A(new_n353_), .B(new_n571_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n571_), .B(new_n635_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n641_), .A2(new_n642_), .A3(G8gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n641_), .B2(G8gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n640_), .B(KEYINPUT40), .C1(new_n643_), .C2(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1325gat));
  NAND3_X1  g448(.A1(new_n634_), .A2(new_n617_), .A3(new_n635_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n650_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT41), .B1(new_n650_), .B2(G15gat), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n623_), .A2(new_n625_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n613_), .A2(G15gat), .ZN(new_n654_));
  OAI22_X1  g453(.A1(new_n651_), .A2(new_n652_), .B1(new_n653_), .B2(new_n654_), .ZN(G1326gat));
  NAND3_X1  g454(.A1(new_n634_), .A2(new_n577_), .A3(new_n635_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(G22gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n656_), .B2(G22gat), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n593_), .A2(G22gat), .ZN(new_n660_));
  OAI22_X1  g459(.A1(new_n658_), .A2(new_n659_), .B1(new_n653_), .B2(new_n660_), .ZN(G1327gat));
  NOR2_X1   g460(.A1(new_n631_), .A2(new_n384_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n347_), .A2(new_n371_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n621_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n666_), .B2(new_n254_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n620_), .A2(new_n619_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT102), .B1(new_n595_), .B2(new_n613_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n418_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT43), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n621_), .A2(new_n672_), .A3(new_n418_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n347_), .A2(new_n371_), .A3(new_n384_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT44), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  INV_X1    g476(.A(new_n675_), .ZN(new_n678_));
  AOI211_X1 g477(.A(new_n677_), .B(new_n678_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n676_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n254_), .A2(G29gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n667_), .B1(new_n680_), .B2(new_n681_), .ZN(G1328gat));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683_));
  INV_X1    g482(.A(G36gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n680_), .B2(new_n571_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n666_), .A2(new_n684_), .A3(new_n571_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT45), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n683_), .B1(new_n685_), .B2(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n676_), .A2(new_n679_), .A3(new_n578_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT46), .B(new_n687_), .C1(new_n690_), .C2(new_n684_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1329gat));
  INV_X1    g491(.A(G43gat), .ZN(new_n693_));
  NOR4_X1   g492(.A1(new_n676_), .A2(new_n679_), .A3(new_n693_), .A4(new_n613_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n665_), .B2(new_n613_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT47), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n680_), .A2(G43gat), .A3(new_n617_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT47), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n695_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1330gat));
  AOI21_X1  g500(.A(G50gat), .B1(new_n666_), .B2(new_n577_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n577_), .A2(G50gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n680_), .B2(new_n703_), .ZN(G1331gat));
  INV_X1    g503(.A(new_n347_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n384_), .A2(new_n371_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n634_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n254_), .A2(G57gat), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(KEYINPUT106), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n708_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n668_), .A2(new_n669_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n371_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n705_), .A2(new_n385_), .A3(new_n418_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(G57gat), .B1(new_n719_), .B2(new_n254_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n711_), .A2(new_n713_), .A3(new_n720_), .ZN(G1332gat));
  OR3_X1    g520(.A1(new_n718_), .A2(G64gat), .A3(new_n578_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G64gat), .B1(new_n708_), .B2(new_n578_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(KEYINPUT48), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(KEYINPUT48), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n724_), .B2(new_n725_), .ZN(G1333gat));
  OR3_X1    g525(.A1(new_n718_), .A2(G71gat), .A3(new_n613_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G71gat), .B1(new_n708_), .B2(new_n613_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(KEYINPUT49), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(KEYINPUT49), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(G1334gat));
  OR3_X1    g530(.A1(new_n718_), .A2(G78gat), .A3(new_n593_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G78gat), .B1(new_n708_), .B2(new_n593_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(KEYINPUT50), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(KEYINPUT50), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n732_), .B1(new_n734_), .B2(new_n735_), .ZN(G1335gat));
  NOR3_X1   g535(.A1(new_n705_), .A2(new_n715_), .A3(new_n384_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n674_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(G85gat), .A3(new_n254_), .ZN(new_n739_));
  NOR4_X1   g538(.A1(new_n714_), .A2(new_n705_), .A3(new_n715_), .A4(new_n663_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n254_), .ZN(new_n741_));
  INV_X1    g540(.A(G85gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(KEYINPUT107), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT107), .B1(new_n741_), .B2(new_n742_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n739_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT108), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n739_), .B(new_n748_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1336gat));
  AOI21_X1  g549(.A(G92gat), .B1(new_n740_), .B2(new_n571_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n571_), .A2(G92gat), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT109), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n751_), .B1(new_n738_), .B2(new_n753_), .ZN(G1337gat));
  NAND3_X1  g553(.A1(new_n740_), .A2(new_n617_), .A3(new_n294_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n738_), .A2(new_n617_), .ZN(new_n756_));
  INV_X1    g555(.A(G99gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT51), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n755_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1338gat));
  NAND3_X1  g561(.A1(new_n740_), .A2(new_n295_), .A3(new_n577_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n674_), .A2(new_n577_), .A3(new_n737_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(G106gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n764_), .B2(G106gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT53), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n770_), .B(new_n763_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1339gat));
  XOR2_X1   g571(.A(new_n706_), .B(KEYINPUT110), .Z(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n343_), .B2(new_n339_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n417_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(new_n417_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n337_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n779_), .A2(new_n371_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n323_), .A2(new_n325_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n303_), .A2(new_n304_), .A3(new_n262_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n320_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n305_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT112), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n328_), .A2(new_n790_), .A3(new_n783_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n326_), .A2(KEYINPUT55), .A3(new_n327_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n306_), .A2(new_n312_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n318_), .B1(new_n793_), .B2(new_n786_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n789_), .A2(new_n791_), .A3(new_n792_), .A4(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n335_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(KEYINPUT56), .A3(new_n335_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n781_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n358_), .A2(new_n360_), .A3(new_n364_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n369_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n363_), .A2(new_n361_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT113), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n802_), .B2(new_n366_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n631_), .B1(new_n800_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n779_), .A2(new_n806_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n795_), .A2(KEYINPUT56), .A3(new_n335_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n335_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n417_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT58), .B(new_n811_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n780_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n807_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(KEYINPUT57), .A3(new_n631_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n810_), .A2(new_n818_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n778_), .B1(new_n823_), .B2(new_n385_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n617_), .A2(new_n618_), .A3(new_n254_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G113gat), .B1(new_n826_), .B2(new_n715_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n814_), .A2(new_n815_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n828_), .A2(new_n418_), .A3(new_n817_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT57), .B1(new_n821_), .B2(new_n631_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT114), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n810_), .A2(new_n818_), .A3(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n822_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n385_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n778_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n825_), .A2(KEYINPUT59), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT59), .B1(new_n824_), .B2(new_n825_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n715_), .A2(G113gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT115), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n827_), .B1(new_n841_), .B2(new_n843_), .ZN(G1340gat));
  NOR2_X1   g643(.A1(new_n705_), .A2(KEYINPUT60), .ZN(new_n845_));
  MUX2_X1   g644(.A(new_n845_), .B(KEYINPUT60), .S(G120gat), .Z(new_n846_));
  NAND2_X1  g645(.A1(new_n826_), .A2(new_n846_), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT116), .Z(new_n848_));
  AOI21_X1  g647(.A(new_n778_), .B1(new_n834_), .B2(new_n385_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n838_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n840_), .B(new_n347_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT117), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G120gat), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n851_), .A2(KEYINPUT117), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n848_), .B1(new_n853_), .B2(new_n854_), .ZN(G1341gat));
  INV_X1    g654(.A(G127gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n826_), .A2(new_n856_), .A3(new_n384_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n839_), .A2(new_n384_), .A3(new_n840_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n859_), .B2(new_n856_), .ZN(G1342gat));
  NAND4_X1  g659(.A1(new_n839_), .A2(G134gat), .A3(new_n418_), .A4(new_n840_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n824_), .A2(new_n631_), .A3(new_n825_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863_));
  OR3_X1    g662(.A1(new_n862_), .A2(new_n863_), .A3(G134gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n862_), .B2(G134gat), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n861_), .A2(new_n864_), .A3(new_n865_), .ZN(G1343gat));
  NAND4_X1  g665(.A1(new_n613_), .A2(new_n578_), .A3(new_n254_), .A4(new_n577_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT119), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n824_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n715_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n347_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g673(.A(new_n870_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT120), .B1(new_n875_), .B2(new_n385_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n870_), .A2(new_n877_), .A3(new_n384_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n879_), .B(new_n881_), .ZN(G1346gat));
  OAI21_X1  g681(.A(G162gat), .B1(new_n875_), .B2(new_n417_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n631_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n870_), .A2(new_n204_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1347gat));
  NOR3_X1   g685(.A1(new_n613_), .A2(new_n578_), .A3(new_n254_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT121), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n593_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n837_), .A2(KEYINPUT125), .A3(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n849_), .B2(new_n889_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n891_), .A2(new_n893_), .A3(new_n491_), .A4(new_n715_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n895_));
  INV_X1    g694(.A(G169gat), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897_));
  INV_X1    g696(.A(new_n888_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n371_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n888_), .A2(KEYINPUT122), .A3(new_n715_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n593_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n896_), .B1(new_n903_), .B2(KEYINPUT123), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n849_), .B2(new_n902_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n895_), .B1(new_n904_), .B2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n577_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n822_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n810_), .A2(new_n818_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(KEYINPUT114), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n384_), .B1(new_n911_), .B2(new_n833_), .ZN(new_n912_));
  OAI211_X1 g711(.A(KEYINPUT123), .B(new_n908_), .C1(new_n912_), .C2(new_n778_), .ZN(new_n913_));
  AND4_X1   g712(.A1(G169gat), .A2(new_n906_), .A3(new_n913_), .A4(new_n895_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n894_), .B1(new_n907_), .B2(new_n914_), .ZN(G1348gat));
  INV_X1    g714(.A(new_n824_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n890_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n917_), .A2(new_n532_), .A3(new_n705_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n891_), .A2(new_n347_), .A3(new_n893_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n532_), .ZN(G1349gat));
  NOR2_X1   g719(.A1(new_n385_), .A2(new_n528_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n891_), .A2(new_n893_), .A3(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n513_), .B1(new_n917_), .B2(new_n385_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n891_), .A2(new_n418_), .A3(new_n893_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(G190gat), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n891_), .A2(new_n893_), .A3(new_n512_), .A4(new_n884_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1351gat));
  NOR3_X1   g727(.A1(new_n617_), .A2(new_n578_), .A3(new_n486_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n824_), .A2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n715_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n932_), .A2(KEYINPUT126), .A3(new_n435_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n931_), .A2(G197gat), .A3(new_n715_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n934_), .A2(KEYINPUT126), .ZN(new_n935_));
  AOI211_X1 g734(.A(new_n933_), .B(new_n935_), .C1(new_n435_), .C2(new_n932_), .ZN(G1352gat));
  NAND2_X1  g735(.A1(new_n931_), .A2(new_n347_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g737(.A1(new_n931_), .A2(new_n384_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT63), .B(G211gat), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT63), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n939_), .A2(new_n942_), .A3(new_n444_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944_));
  OR2_X1    g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n944_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n941_), .B1(new_n945_), .B2(new_n946_), .ZN(G1354gat));
  INV_X1    g746(.A(new_n931_), .ZN(new_n948_));
  OAI21_X1  g747(.A(G218gat), .B1(new_n948_), .B2(new_n417_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n931_), .A2(new_n442_), .A3(new_n884_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1355gat));
endmodule


