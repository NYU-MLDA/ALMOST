//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n919_, new_n921_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_;
  XNOR2_X1  g000(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G190gat), .B(G218gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT75), .ZN(new_n205_));
  XOR2_X1   g004(.A(G134gat), .B(G162gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT36), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR3_X1   g012(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n210_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  INV_X1    g015(.A(G99gat), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n219_), .A2(KEYINPUT66), .A3(new_n212_), .A4(new_n211_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n221_), .A2(KEYINPUT67), .A3(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(G85gat), .B(G92gat), .Z(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n228_), .B1(new_n215_), .B2(new_n220_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(KEYINPUT67), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT68), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n233_), .B1(new_n236_), .B2(KEYINPUT67), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n215_), .A2(new_n220_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(new_n228_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n231_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n227_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n226_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n223_), .A2(new_n225_), .A3(KEYINPUT69), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n246_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n245_), .B1(new_n250_), .B2(new_n221_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT70), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT8), .B1(new_n251_), .B2(KEYINPUT70), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n238_), .B(new_n244_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G29gat), .B(G36gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G43gat), .B(G50gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n223_), .A2(new_n225_), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT10), .B(G99gat), .Z(new_n260_));
  AOI21_X1  g059(.A(new_n259_), .B1(new_n218_), .B2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT64), .B1(G85gat), .B2(G92gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT9), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n263_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n264_), .B(new_n265_), .C1(G85gat), .C2(G92gat), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n255_), .A2(new_n258_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n255_), .A2(KEYINPUT73), .A3(new_n258_), .A4(new_n268_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G232gat), .A2(G233gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT34), .Z(new_n274_));
  INV_X1    g073(.A(KEYINPUT35), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT74), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n271_), .A2(KEYINPUT74), .A3(new_n272_), .A4(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n255_), .A2(new_n268_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n258_), .B(KEYINPUT15), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT72), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n279_), .A2(new_n280_), .A3(new_n285_), .A4(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n274_), .A2(new_n275_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n277_), .A2(new_n289_), .A3(new_n286_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n209_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n207_), .A2(new_n208_), .ZN(new_n294_));
  AOI211_X1 g093(.A(new_n291_), .B(new_n294_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n203_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n294_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n290_), .A2(new_n292_), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n291_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n298_), .B(new_n202_), .C1(new_n299_), .C2(new_n209_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G127gat), .B(G155gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT16), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G183gat), .B(G211gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT17), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G15gat), .B(G22gat), .ZN(new_n308_));
  INV_X1    g107(.A(G1gat), .ZN(new_n309_));
  INV_X1    g108(.A(G8gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT14), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G1gat), .B(G8gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G231gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G57gat), .B(G64gat), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n317_), .A2(KEYINPUT11), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(KEYINPUT11), .ZN(new_n319_));
  XOR2_X1   g118(.A(G71gat), .B(G78gat), .Z(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n319_), .A2(new_n320_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n316_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n307_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n327_), .B1(new_n326_), .B2(new_n325_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n306_), .A2(KEYINPUT17), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n329_), .B(KEYINPUT77), .Z(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n325_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n302_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n323_), .B(new_n326_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n255_), .A2(new_n268_), .A3(new_n334_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n223_), .A2(new_n225_), .A3(KEYINPUT69), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT69), .B1(new_n223_), .B2(new_n225_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n227_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n231_), .B1(new_n241_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n232_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n239_), .A2(new_n242_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n341_), .A2(new_n252_), .B1(new_n342_), .B2(KEYINPUT68), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n267_), .B1(new_n343_), .B2(new_n244_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n324_), .A2(KEYINPUT12), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n335_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n334_), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT12), .B1(new_n281_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G230gat), .A2(G233gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n346_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n281_), .A2(new_n347_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n349_), .B1(new_n352_), .B2(new_n335_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G120gat), .B(G148gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT5), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G176gat), .B(G204gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  OR3_X1    g156(.A1(new_n351_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT13), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(KEYINPUT13), .A3(new_n359_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n314_), .B(new_n258_), .Z(new_n365_));
  NAND2_X1  g164(.A1(G229gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT78), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n282_), .A2(new_n314_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n314_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n258_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n372_), .A3(new_n366_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G113gat), .B(G141gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G169gat), .B(G197gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n377_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n364_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT99), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT96), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT20), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT23), .ZN(new_n394_));
  INV_X1    g193(.A(G169gat), .ZN(new_n395_));
  INV_X1    g194(.A(G176gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n397_), .A2(KEYINPUT24), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G169gat), .A2(G176gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(KEYINPUT24), .A3(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n394_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT26), .B(G190gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT25), .B(G183gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n394_), .B1(G183gat), .B2(G190gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT81), .B(G176gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT22), .B(G169gat), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n406_), .A2(new_n407_), .B1(G169gat), .B2(G176gat), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n401_), .A2(new_n404_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT89), .ZN(new_n410_));
  INV_X1    g209(.A(G197gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(G204gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(G204gat), .ZN(new_n413_));
  INV_X1    g212(.A(G204gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n412_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n416_), .A2(KEYINPUT21), .ZN(new_n417_));
  XOR2_X1   g216(.A(G211gat), .B(G218gat), .Z(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(G197gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n413_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(KEYINPUT21), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G211gat), .B(G218gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT21), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n417_), .A2(new_n421_), .B1(new_n416_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n392_), .B1(new_n409_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT98), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT94), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT26), .B(G190gat), .Z(new_n429_));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT80), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT26), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT79), .B1(new_n433_), .B2(G190gat), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n431_), .A2(new_n432_), .A3(new_n434_), .A4(new_n403_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n434_), .B(new_n403_), .C1(new_n402_), .C2(KEYINPUT79), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT80), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n437_), .A3(new_n401_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n405_), .A2(new_n408_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT82), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n442_), .A3(new_n439_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n420_), .A2(KEYINPUT21), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n445_), .B(new_n422_), .C1(new_n416_), .C2(KEYINPUT21), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n424_), .A2(new_n416_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n428_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n438_), .A2(new_n442_), .A3(new_n439_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n442_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n428_), .B(new_n448_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n427_), .B1(new_n449_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G226gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT19), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n401_), .A2(new_n404_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n439_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(KEYINPUT93), .A3(new_n448_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT93), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n409_), .B2(new_n425_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n392_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n441_), .A2(new_n443_), .A3(new_n425_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n456_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n391_), .B1(new_n457_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n426_), .A2(new_n465_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n449_), .B2(new_n453_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n465_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n472_), .A3(new_n391_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G85gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT0), .B(G57gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G127gat), .B(G134gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G113gat), .B(G120gat), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n479_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT84), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT3), .ZN(new_n485_));
  INV_X1    g284(.A(G141gat), .ZN(new_n486_));
  INV_X1    g285(.A(G148gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G141gat), .A2(G148gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT2), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n488_), .A2(new_n491_), .A3(new_n492_), .A4(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(G155gat), .A2(G162gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G155gat), .A2(G162gat), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(KEYINPUT1), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT1), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(G155gat), .A3(G162gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n501_), .A3(new_n495_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n486_), .A2(new_n487_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n489_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n480_), .A2(KEYINPUT84), .A3(new_n481_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n484_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n498_), .A2(new_n504_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n482_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G225gat), .A2(G233gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n513_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n477_), .B(new_n512_), .C1(new_n517_), .C2(new_n511_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n477_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n515_), .A2(new_n516_), .A3(new_n511_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n512_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n473_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n383_), .B1(new_n467_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT98), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n426_), .B(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n448_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT94), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(new_n529_), .B2(new_n452_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n466_), .B1(new_n530_), .B2(new_n465_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n391_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n533_), .A2(KEYINPUT99), .A3(new_n523_), .A4(new_n473_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n477_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(new_n517_), .B2(new_n511_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n522_), .A2(KEYINPUT97), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(KEYINPUT33), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n470_), .A2(new_n472_), .A3(new_n390_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n468_), .B1(new_n529_), .B2(new_n452_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n389_), .B1(new_n540_), .B2(new_n471_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT33), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n522_), .A2(KEYINPUT97), .A3(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .A4(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n525_), .A2(new_n534_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT28), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n508_), .B2(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n505_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G22gat), .B(G50gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n548_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G78gat), .B(G106gat), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT90), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n547_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n425_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n558_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(KEYINPUT90), .A3(new_n448_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT87), .B(G228gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT88), .B(G233gat), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n561_), .A3(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n560_), .A2(new_n448_), .A3(KEYINPUT90), .A4(new_n564_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n554_), .B1(new_n556_), .B2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n556_), .B1(new_n568_), .B2(KEYINPUT91), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT91), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n566_), .A2(new_n571_), .A3(new_n567_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n570_), .A2(KEYINPUT92), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT92), .B1(new_n570_), .B2(new_n572_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n569_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n554_), .A2(KEYINPUT86), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n554_), .A2(KEYINPUT86), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n568_), .A2(new_n556_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n566_), .A2(new_n555_), .A3(new_n567_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT83), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT30), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n450_), .A2(new_n451_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT30), .B1(new_n441_), .B2(new_n443_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n583_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n584_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n441_), .A2(KEYINPUT30), .A3(new_n443_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT83), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G71gat), .B(G99gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(G43gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G227gat), .A2(G233gat), .ZN(new_n593_));
  INV_X1    g392(.A(G15gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n592_), .B(new_n595_), .Z(new_n596_));
  NAND3_X1  g395(.A1(new_n587_), .A2(new_n590_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n484_), .A2(new_n506_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n598_), .A2(KEYINPUT31), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(KEYINPUT31), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n599_), .A2(KEYINPUT85), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(KEYINPUT83), .B1(new_n588_), .B2(new_n589_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n596_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n600_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT85), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n597_), .A2(new_n604_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n597_), .B2(new_n604_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n575_), .B(new_n582_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n545_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n569_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n570_), .A2(new_n572_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT92), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n570_), .A2(KEYINPUT92), .A3(new_n572_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n582_), .ZN(new_n620_));
  OAI22_X1  g419(.A1(new_n619_), .A2(new_n620_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n597_), .A2(new_n604_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n607_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n597_), .A2(new_n604_), .A3(new_n608_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n575_), .A2(new_n623_), .A3(new_n624_), .A4(new_n582_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n466_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n627_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT27), .B(new_n539_), .C1(new_n628_), .C2(new_n390_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT27), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n390_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n540_), .A2(new_n389_), .A3(new_n471_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n523_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n629_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n626_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n613_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n382_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n333_), .A2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT100), .Z(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n309_), .A3(new_n523_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(KEYINPUT105), .A2(KEYINPUT38), .ZN(new_n642_));
  AND2_X1   g441(.A1(KEYINPUT105), .A2(KEYINPUT38), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT101), .B1(new_n293_), .B2(new_n295_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n298_), .B(new_n646_), .C1(new_n299_), .C2(new_n209_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n637_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT102), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n651_), .A3(new_n637_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n332_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT103), .B1(new_n653_), .B2(new_n382_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(KEYINPUT103), .A3(new_n382_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n523_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n658_), .A2(KEYINPUT104), .A3(G1gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT104), .B1(new_n658_), .B2(G1gat), .ZN(new_n660_));
  OAI221_X1 g459(.A(new_n644_), .B1(new_n642_), .B2(new_n641_), .C1(new_n659_), .C2(new_n660_), .ZN(G1324gat));
  NAND2_X1  g460(.A1(new_n629_), .A2(new_n633_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n640_), .A2(new_n310_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n650_), .A2(new_n652_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n332_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n664_), .A2(new_n382_), .A3(new_n665_), .A4(new_n662_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n666_), .A2(KEYINPUT106), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n310_), .B1(new_n666_), .B2(KEYINPUT106), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n663_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(G1325gat));
  NOR2_X1   g473(.A1(new_n609_), .A2(new_n610_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n640_), .A2(new_n594_), .A3(new_n675_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n653_), .A2(KEYINPUT103), .A3(new_n382_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n677_), .B2(new_n654_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n678_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(new_n678_), .B2(G15gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT107), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n683_), .B(new_n676_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1326gat));
  INV_X1    g484(.A(G22gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n619_), .A2(new_n620_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n640_), .A2(new_n686_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n657_), .A2(new_n688_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(G22gat), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT42), .B(new_n686_), .C1(new_n657_), .C2(new_n688_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(G1327gat));
  NAND3_X1  g493(.A1(new_n296_), .A2(new_n300_), .A3(new_n637_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT43), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n296_), .A2(new_n300_), .A3(new_n637_), .A4(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n364_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(new_n380_), .A3(new_n332_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT44), .B1(new_n699_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n704_), .B(new_n701_), .C1(new_n696_), .C2(new_n698_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n703_), .A2(new_n705_), .A3(new_n634_), .ZN(new_n706_));
  INV_X1    g505(.A(G29gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n648_), .A2(new_n665_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n638_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n708_), .A2(KEYINPUT108), .A3(new_n638_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n523_), .A2(new_n707_), .ZN(new_n714_));
  OAI22_X1  g513(.A1(new_n706_), .A2(new_n707_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716_));
  INV_X1    g515(.A(new_n662_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n703_), .A2(new_n705_), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719_));
  OAI21_X1  g518(.A(G36gat), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n699_), .A2(new_n702_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n704_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n699_), .A2(KEYINPUT44), .A3(new_n702_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n662_), .A3(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(KEYINPUT109), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n716_), .B1(new_n720_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n718_), .A2(new_n719_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(KEYINPUT109), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(KEYINPUT110), .A4(G36gat), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n717_), .A2(G36gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n711_), .A2(new_n712_), .A3(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n726_), .A2(new_n729_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n727_), .A2(new_n728_), .A3(G36gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n733_), .B1(new_n741_), .B2(new_n716_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n742_), .A2(new_n736_), .A3(new_n737_), .A4(new_n729_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n740_), .A2(new_n743_), .ZN(G1329gat));
  NOR4_X1   g543(.A1(new_n713_), .A2(G43gat), .A3(new_n610_), .A4(new_n609_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n722_), .A2(new_n675_), .A3(new_n723_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(G43gat), .B2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g547(.A1(new_n703_), .A2(new_n705_), .A3(new_n687_), .ZN(new_n749_));
  INV_X1    g548(.A(G50gat), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n687_), .A2(G50gat), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT113), .ZN(new_n752_));
  OAI22_X1  g551(.A1(new_n749_), .A2(new_n750_), .B1(new_n713_), .B2(new_n752_), .ZN(G1331gat));
  NOR2_X1   g552(.A1(new_n700_), .A2(new_n380_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n653_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(G57gat), .A3(new_n523_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(KEYINPUT114), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(KEYINPUT114), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n754_), .A2(new_n637_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n333_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n523_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n757_), .A2(new_n758_), .A3(new_n762_), .ZN(G1332gat));
  INV_X1    g562(.A(G64gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n755_), .B2(new_n662_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT48), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n761_), .A2(new_n764_), .A3(new_n662_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1333gat));
  NAND2_X1  g567(.A1(new_n755_), .A2(new_n675_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G71gat), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n609_), .A2(new_n610_), .A3(G71gat), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT116), .Z(new_n774_));
  OAI21_X1  g573(.A(new_n772_), .B1(new_n760_), .B2(new_n774_), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n755_), .A2(new_n688_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G78gat), .ZN(new_n777_));
  XNOR2_X1  g576(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n777_), .B(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n687_), .A2(G78gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n760_), .B2(new_n780_), .ZN(G1335gat));
  AND2_X1   g580(.A1(new_n759_), .A2(new_n708_), .ZN(new_n782_));
  INV_X1    g581(.A(G85gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n523_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n699_), .A2(new_n332_), .A3(new_n754_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n523_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n786_), .B2(new_n783_), .ZN(G1336gat));
  INV_X1    g586(.A(G92gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n782_), .A2(new_n788_), .A3(new_n662_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n785_), .A2(new_n662_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(new_n788_), .ZN(G1337gat));
  AOI21_X1  g590(.A(new_n217_), .B1(new_n785_), .B2(new_n675_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT118), .ZN(new_n793_));
  NAND2_X1  g592(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n782_), .A2(new_n260_), .A3(new_n675_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n796_), .B(new_n797_), .Z(G1338gat));
  AOI21_X1  g597(.A(new_n218_), .B1(new_n785_), .B2(new_n688_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT52), .Z(new_n800_));
  NAND3_X1  g599(.A1(new_n782_), .A2(new_n218_), .A3(new_n688_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g602(.A(new_n625_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n662_), .A2(new_n634_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n365_), .A2(new_n366_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n370_), .A2(new_n372_), .A3(new_n367_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n377_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n378_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n360_), .A2(new_n809_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n255_), .A2(new_n268_), .A3(new_n334_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n345_), .B1(new_n255_), .B2(new_n268_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT12), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n344_), .B2(new_n334_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n349_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n349_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n350_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n351_), .A2(new_n820_), .A3(KEYINPUT55), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT56), .B1(new_n822_), .B2(new_n357_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824_));
  INV_X1    g623(.A(new_n357_), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n824_), .B(new_n825_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n823_), .A2(new_n826_), .A3(KEYINPUT121), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n351_), .B1(KEYINPUT55), .B2(new_n820_), .ZN(new_n828_));
  NOR4_X1   g627(.A1(new_n346_), .A2(new_n348_), .A3(new_n818_), .A4(new_n350_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n357_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(KEYINPUT121), .A3(new_n824_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n358_), .A2(new_n380_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n810_), .B1(new_n827_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n648_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n830_), .A2(new_n824_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n822_), .A2(KEYINPUT56), .A3(new_n357_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n809_), .A2(new_n358_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT58), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n843_), .B(new_n840_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n835_), .A2(new_n836_), .B1(new_n845_), .B2(new_n302_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n834_), .A2(KEYINPUT57), .A3(new_n648_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n665_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n381_), .A2(new_n665_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT120), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n301_), .A2(new_n700_), .A3(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT54), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n804_), .B(new_n805_), .C1(new_n848_), .C2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(G113gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n380_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n858_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n831_), .A2(new_n832_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n837_), .A2(new_n861_), .A3(new_n838_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n860_), .A2(new_n862_), .B1(new_n360_), .B2(new_n809_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n645_), .A2(new_n647_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n836_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n845_), .A2(new_n302_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n847_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n332_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n852_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n869_), .A2(KEYINPUT59), .A3(new_n804_), .A4(new_n805_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n381_), .B1(new_n859_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n857_), .B1(new_n871_), .B2(new_n856_), .ZN(G1340gat));
  AOI21_X1  g671(.A(new_n700_), .B1(new_n859_), .B2(new_n870_), .ZN(new_n873_));
  INV_X1    g672(.A(G120gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(KEYINPUT60), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n700_), .B2(KEYINPUT60), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n877_), .B2(new_n876_), .ZN(new_n879_));
  OAI22_X1  g678(.A1(new_n873_), .A2(new_n874_), .B1(new_n854_), .B2(new_n879_), .ZN(G1341gat));
  INV_X1    g679(.A(G127gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n855_), .A2(new_n881_), .A3(new_n665_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n332_), .B1(new_n859_), .B2(new_n870_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT123), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n886_), .B(new_n882_), .C1(new_n883_), .C2(new_n881_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1342gat));
  INV_X1    g687(.A(G134gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n855_), .A2(new_n889_), .A3(new_n864_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n301_), .B1(new_n859_), .B2(new_n870_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1343gat));
  AOI21_X1  g691(.A(new_n621_), .B1(new_n868_), .B2(new_n852_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n805_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n381_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n486_), .ZN(G1344gat));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n700_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n487_), .ZN(G1345gat));
  INV_X1    g697(.A(new_n621_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n869_), .A2(new_n665_), .A3(new_n899_), .A4(new_n805_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT124), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT61), .B(G155gat), .Z(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  OAI21_X1  g702(.A(G162gat), .B1(new_n894_), .B2(new_n301_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n648_), .A2(G162gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n894_), .B2(new_n905_), .ZN(G1347gat));
  AOI21_X1  g705(.A(new_n625_), .B1(new_n868_), .B2(new_n852_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n717_), .A2(new_n523_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n381_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n911_));
  OR3_X1    g710(.A1(new_n910_), .A2(new_n395_), .A3(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n910_), .B2(new_n395_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n407_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(G1348gat));
  NAND3_X1  g714(.A1(new_n907_), .A2(new_n364_), .A3(new_n908_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n396_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n406_), .B2(new_n916_), .ZN(G1349gat));
  NOR2_X1   g717(.A1(new_n909_), .A2(new_n332_), .ZN(new_n919_));
  MUX2_X1   g718(.A(G183gat), .B(new_n403_), .S(new_n919_), .Z(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n909_), .B2(new_n301_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n864_), .A2(new_n402_), .ZN(new_n922_));
  XOR2_X1   g721(.A(new_n922_), .B(KEYINPUT126), .Z(new_n923_));
  OAI21_X1  g722(.A(new_n921_), .B1(new_n909_), .B2(new_n923_), .ZN(G1351gat));
  NAND2_X1  g723(.A1(new_n893_), .A2(new_n908_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n381_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(new_n411_), .ZN(G1352gat));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n700_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(new_n414_), .ZN(G1353gat));
  INV_X1    g728(.A(new_n925_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT63), .B(G211gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n930_), .A2(new_n665_), .A3(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933_));
  OAI22_X1  g732(.A1(new_n925_), .A2(new_n332_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n933_), .B1(new_n932_), .B2(new_n934_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1354gat));
  OR3_X1    g736(.A1(new_n925_), .A2(G218gat), .A3(new_n648_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G218gat), .B1(new_n925_), .B2(new_n301_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1355gat));
endmodule


