//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n967_, new_n968_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n989_, new_n990_, new_n991_, new_n992_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_;
  XNOR2_X1  g000(.A(KEYINPUT79), .B(KEYINPUT28), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G22gat), .B(G50gat), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G141gat), .ZN(new_n206_));
  INV_X1    g005(.A(G148gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n208_), .A2(KEYINPUT3), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT77), .B1(new_n208_), .B2(KEYINPUT3), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .A4(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G155gat), .B(G162gat), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n210_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n208_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n214_), .A2(KEYINPUT76), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n222_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n219_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n220_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT78), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n218_), .A2(new_n219_), .B1(new_n228_), .B2(new_n226_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n205_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  AOI211_X1 g036(.A(KEYINPUT29), .B(new_n204_), .C1(new_n231_), .C2(new_n234_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n203_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n230_), .A2(KEYINPUT78), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n232_), .A2(new_n233_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n236_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n204_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n235_), .A2(new_n236_), .A3(new_n205_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n202_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n239_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n231_), .A2(KEYINPUT29), .A3(new_n234_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G197gat), .B(G204gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(G197gat), .A2(G204gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G197gat), .A2(G204gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(KEYINPUT21), .A3(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n255_), .A2(new_n256_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n258_), .A3(KEYINPUT82), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(G233gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT81), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n265_), .A2(G228gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(G228gat), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n264_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n263_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n249_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n259_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(KEYINPUT83), .A3(new_n269_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT83), .B1(new_n272_), .B2(new_n269_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n271_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G78gat), .B(G106gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n271_), .B(new_n279_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n248_), .A2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n239_), .A2(new_n245_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT80), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n286_));
  INV_X1    g085(.A(new_n259_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n230_), .B2(KEYINPUT29), .ZN(new_n288_));
  INV_X1    g087(.A(new_n269_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n286_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n290_), .A2(new_n273_), .B1(new_n249_), .B2(new_n270_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT84), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n277_), .B1(new_n291_), .B2(KEYINPUT84), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n283_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n280_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n291_), .A2(KEYINPUT85), .A3(new_n279_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n295_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT84), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n279_), .B1(new_n276_), .B2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n246_), .B1(new_n303_), .B2(new_n292_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n297_), .A2(new_n298_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT86), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n285_), .B1(new_n301_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT95), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT19), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT87), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n257_), .A2(new_n258_), .A3(KEYINPUT82), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT82), .B1(new_n257_), .B2(new_n258_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G183gat), .ZN(new_n315_));
  INV_X1    g114(.A(G190gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT23), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G183gat), .A3(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n316_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n320_), .A2(new_n321_), .B1(G169gat), .B2(G176gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT22), .B(G169gat), .ZN(new_n323_));
  INV_X1    g122(.A(G176gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT73), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n323_), .A2(new_n327_), .A3(new_n324_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n322_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n317_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n319_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n319_), .A2(new_n331_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n330_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT25), .B(G183gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT26), .B(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(KEYINPUT24), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT24), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n337_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n329_), .B1(new_n334_), .B2(new_n344_), .ZN(new_n345_));
  OAI211_X1 g144(.A(KEYINPUT88), .B(KEYINPUT20), .C1(new_n314_), .C2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n337_), .A2(new_n341_), .A3(new_n343_), .A4(new_n320_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT89), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n335_), .A2(new_n336_), .B1(new_n342_), .B2(new_n338_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n350_), .A2(KEYINPUT89), .A3(new_n341_), .A4(new_n320_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n321_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n340_), .B(new_n325_), .C1(new_n334_), .C2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n259_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n346_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n332_), .A2(new_n333_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n317_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n341_), .A3(new_n350_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(new_n329_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT88), .B1(new_n361_), .B2(KEYINPUT20), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n311_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n314_), .A2(new_n345_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n310_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n352_), .A2(new_n287_), .A3(new_n354_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n368_), .A2(KEYINPUT20), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n363_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT27), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n346_), .A2(new_n356_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n311_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n362_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n325_), .A2(new_n340_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n359_), .B2(new_n321_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n347_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n380_));
  OAI211_X1 g179(.A(KEYINPUT94), .B(KEYINPUT20), .C1(new_n379_), .C2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n368_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n354_), .A2(new_n287_), .A3(new_n347_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT94), .B1(new_n383_), .B2(KEYINPUT20), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n310_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n367_), .B1(new_n377_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n308_), .B1(new_n373_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n367_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n357_), .A2(new_n311_), .A3(new_n362_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n369_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n393_), .A2(KEYINPUT95), .A3(KEYINPUT27), .A4(new_n372_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT27), .ZN(new_n395_));
  INV_X1    g194(.A(new_n372_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n367_), .B1(new_n363_), .B2(new_n371_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n389_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G127gat), .B(G134gat), .Z(new_n400_));
  XOR2_X1   g199(.A(G113gat), .B(G120gat), .Z(new_n401_));
  XOR2_X1   g200(.A(new_n400_), .B(new_n401_), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT74), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT30), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT31), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408_));
  INV_X1    g207(.A(G71gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G99gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n345_), .B(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT75), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n407_), .A2(new_n412_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n403_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n415_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT75), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n402_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n231_), .A2(new_n234_), .A3(new_n402_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n403_), .A2(new_n232_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(KEYINPUT4), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT90), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n424_), .A2(new_n428_), .A3(KEYINPUT4), .A4(new_n425_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G225gat), .A2(G233gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n431_), .B(KEYINPUT91), .Z(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(new_n424_), .B2(KEYINPUT4), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G1gat), .B(G29gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G57gat), .B(G85gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n424_), .A2(new_n425_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n440_), .B1(new_n441_), .B2(new_n432_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n435_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n440_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n433_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n441_), .A2(new_n432_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n423_), .A2(new_n450_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n307_), .A2(new_n399_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n363_), .A2(new_n371_), .A3(new_n453_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n442_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT93), .B1(new_n459_), .B2(KEYINPUT33), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT93), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n461_), .B(new_n462_), .C1(new_n446_), .C2(new_n442_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n446_), .A2(new_n462_), .A3(new_n442_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n432_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n445_), .B1(new_n441_), .B2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n424_), .A2(KEYINPUT4), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(new_n432_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n430_), .B2(new_n469_), .ZN(new_n470_));
  NOR4_X1   g269(.A1(new_n465_), .A2(new_n396_), .A3(new_n470_), .A4(new_n397_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n458_), .B1(new_n464_), .B2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n300_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n304_), .A2(KEYINPUT86), .A3(new_n305_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n473_), .A2(new_n474_), .B1(new_n284_), .B2(new_n282_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n423_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n450_), .A2(new_n389_), .A3(new_n394_), .A4(new_n398_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n307_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n452_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT69), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT70), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G1gat), .B(G8gat), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G29gat), .B(G36gat), .Z(new_n491_));
  XOR2_X1   g290(.A(G43gat), .B(G50gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n482_), .A2(new_n488_), .A3(new_n486_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n493_), .B(KEYINPUT15), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n490_), .A2(new_n494_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n495_), .B(new_n496_), .C1(new_n498_), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n496_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n495_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n493_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n501_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n479_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G127gat), .B(G155gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT16), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G183gat), .B(G211gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT71), .ZN(new_n522_));
  AND2_X1   g321(.A1(G231gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n499_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G57gat), .B(G64gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G71gat), .B(G78gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(KEYINPUT11), .ZN(new_n527_));
  XOR2_X1   g326(.A(G71gat), .B(G78gat), .Z(new_n528_));
  INV_X1    g327(.A(G64gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(G57gat), .ZN(new_n530_));
  INV_X1    g329(.A(G57gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(G64gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n532_), .A3(KEYINPUT11), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n525_), .A2(KEYINPUT11), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n527_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT65), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT65), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n538_), .B(new_n527_), .C1(new_n534_), .C2(new_n535_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n524_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n524_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n530_), .A2(new_n532_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT11), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(new_n533_), .A3(new_n528_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n538_), .B1(new_n547_), .B2(new_n527_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n542_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n522_), .A2(new_n541_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n542_), .A2(new_n536_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n519_), .A2(new_n520_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n524_), .A2(new_n527_), .A3(new_n547_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(G85gat), .ZN(new_n557_));
  INV_X1    g356(.A(G92gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G85gat), .A2(G92gat), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  OR3_X1    g360(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(G99gat), .B2(G106gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(KEYINPUT6), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n562_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT64), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT64), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n561_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT8), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n565_), .A2(KEYINPUT6), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n563_), .A2(G99gat), .A3(G106gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n578_), .A2(new_n562_), .A3(new_n570_), .A4(new_n571_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(KEYINPUT8), .A3(new_n561_), .ZN(new_n580_));
  OR2_X1    g379(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n581_));
  INV_X1    g380(.A(G106gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n559_), .A2(KEYINPUT9), .A3(new_n560_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n560_), .A2(KEYINPUT9), .ZN(new_n586_));
  AND4_X1   g385(.A1(new_n578_), .A2(new_n584_), .A3(new_n585_), .A4(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n575_), .A2(new_n580_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n497_), .A2(new_n589_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n579_), .A2(KEYINPUT8), .A3(new_n561_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT8), .B1(new_n579_), .B2(new_n561_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n591_), .A2(new_n592_), .A3(new_n587_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n493_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT34), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n590_), .A2(new_n594_), .A3(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(KEYINPUT35), .A3(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n590_), .A2(new_n600_), .A3(new_n594_), .A4(new_n597_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n599_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n599_), .A2(new_n601_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n604_), .B(KEYINPUT36), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n606_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT37), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n612_), .B(new_n606_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n556_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n593_), .A2(new_n540_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n549_), .A2(new_n589_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT66), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n619_), .B(new_n621_), .C1(new_n618_), .C2(new_n617_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT67), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n547_), .A2(KEYINPUT12), .A3(new_n527_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n593_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n624_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n589_), .A2(KEYINPUT67), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT12), .B1(new_n549_), .B2(new_n589_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n617_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(new_n630_), .A3(new_n620_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n622_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT5), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n634_), .B(new_n635_), .Z(new_n636_));
  NAND2_X1  g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n636_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n622_), .A2(new_n631_), .A3(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(KEYINPUT68), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT68), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n632_), .A2(new_n641_), .A3(new_n636_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n640_), .A2(KEYINPUT13), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT13), .B1(new_n640_), .B2(new_n642_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n615_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n515_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  AOI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(KEYINPUT96), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n449_), .A3(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(KEYINPUT96), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n645_), .A2(new_n514_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n556_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n610_), .B(KEYINPUT97), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT98), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT99), .B1(new_n479_), .B2(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n389_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n475_), .A2(new_n661_), .A3(new_n450_), .A4(new_n423_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n418_), .A2(new_n422_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n455_), .A2(new_n456_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n449_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n460_), .A2(new_n463_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n435_), .A2(KEYINPUT33), .A3(new_n443_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n430_), .A2(new_n469_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n467_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n363_), .A2(new_n371_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n390_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n667_), .A2(new_n670_), .A3(new_n372_), .A4(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n665_), .B1(new_n666_), .B2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n663_), .B1(new_n307_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n473_), .A2(new_n474_), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n661_), .A2(new_n450_), .B1(new_n676_), .B2(new_n285_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n662_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n658_), .B(KEYINPUT98), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n657_), .B1(new_n660_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n449_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n683_), .A2(KEYINPUT100), .A3(G1gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT100), .B1(new_n683_), .B2(G1gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n653_), .B1(new_n684_), .B2(new_n685_), .ZN(G1324gat));
  AND3_X1   g485(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n679_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n399_), .B(new_n656_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G8gat), .B1(new_n689_), .B2(KEYINPUT101), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n682_), .B2(new_n399_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT39), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n682_), .A2(new_n691_), .A3(new_n399_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(KEYINPUT101), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT39), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .A4(G8gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n693_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n648_), .A2(new_n484_), .A3(new_n399_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT40), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n698_), .A2(KEYINPUT40), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1325gat));
  OR3_X1    g503(.A1(new_n647_), .A2(G15gat), .A3(new_n663_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n682_), .A2(new_n423_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n706_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT41), .B1(new_n706_), .B2(G15gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(G1326gat));
  OR3_X1    g508(.A1(new_n647_), .A2(G22gat), .A3(new_n475_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n682_), .A2(new_n307_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G22gat), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(KEYINPUT42), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(KEYINPUT42), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(G1327gat));
  NAND2_X1  g514(.A1(new_n658_), .A2(new_n556_), .ZN(new_n716_));
  NOR4_X1   g515(.A1(new_n479_), .A2(new_n514_), .A3(new_n645_), .A4(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G29gat), .B1(new_n717_), .B2(new_n449_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n611_), .A2(new_n613_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n719_), .B2(KEYINPUT102), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n396_), .A2(new_n470_), .A3(new_n397_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n722_), .A2(new_n667_), .A3(new_n460_), .A4(new_n463_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n475_), .A2(new_n665_), .A3(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n478_), .A3(new_n663_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n719_), .B(new_n721_), .C1(new_n725_), .C2(new_n662_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n719_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n720_), .B1(new_n678_), .B2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n556_), .B(new_n654_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT103), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n729_), .A2(new_n731_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n449_), .A2(G29gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n718_), .B1(new_n734_), .B2(new_n735_), .ZN(G1328gat));
  INV_X1    g535(.A(G36gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n717_), .A2(new_n737_), .A3(new_n399_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT45), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n661_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(new_n737_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT46), .B(new_n739_), .C1(new_n740_), .C2(new_n737_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1329gat));
  INV_X1    g544(.A(G43gat), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n663_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n717_), .A2(new_n423_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT104), .B1(new_n750_), .B2(new_n746_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT104), .B(new_n748_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT47), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n749_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n756_), .B(new_n757_), .C1(new_n749_), .C2(new_n751_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(new_n758_), .ZN(G1330gat));
  AOI21_X1  g558(.A(G50gat), .B1(new_n717_), .B2(new_n307_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n307_), .A2(G50gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n734_), .B2(new_n761_), .ZN(G1331gat));
  NAND2_X1  g561(.A1(new_n678_), .A2(new_n514_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n763_), .A2(KEYINPUT105), .ZN(new_n764_));
  INV_X1    g563(.A(new_n645_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n763_), .B2(KEYINPUT105), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(new_n615_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G57gat), .B1(new_n768_), .B2(new_n449_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n645_), .A2(new_n514_), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n556_), .B(new_n770_), .C1(new_n660_), .C2(new_n681_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n531_), .B1(new_n449_), .B2(KEYINPUT106), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(KEYINPUT106), .B2(new_n531_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n769_), .B1(new_n771_), .B2(new_n773_), .ZN(G1332gat));
  NAND3_X1  g573(.A1(new_n768_), .A2(new_n529_), .A3(new_n399_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n771_), .A2(new_n399_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G64gat), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT48), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(KEYINPUT48), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1333gat));
  NAND3_X1  g579(.A1(new_n768_), .A2(new_n409_), .A3(new_n423_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n771_), .A2(new_n423_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G71gat), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(KEYINPUT49), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT49), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1334gat));
  INV_X1    g585(.A(G78gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n768_), .A2(new_n787_), .A3(new_n307_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n771_), .A2(new_n307_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(G78gat), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n790_), .A2(KEYINPUT50), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(KEYINPUT50), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(G1335gat));
  INV_X1    g592(.A(new_n716_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n764_), .A2(new_n766_), .A3(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n557_), .B1(new_n795_), .B2(new_n450_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT107), .Z(new_n797_));
  OR2_X1    g596(.A1(new_n726_), .A2(new_n728_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n556_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n770_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n801_), .A2(new_n557_), .A3(new_n450_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n797_), .A2(new_n802_), .ZN(G1336gat));
  INV_X1    g602(.A(new_n795_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G92gat), .B1(new_n804_), .B2(new_n399_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n801_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n399_), .A2(G92gat), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT108), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n805_), .B1(new_n806_), .B2(new_n808_), .ZN(G1337gat));
  OAI21_X1  g608(.A(G99gat), .B1(new_n801_), .B2(new_n663_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n423_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n804_), .A2(KEYINPUT109), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT109), .B1(new_n804_), .B2(new_n812_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT51), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n817_), .B(new_n810_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1338gat));
  XNOR2_X1  g618(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n307_), .B(new_n800_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G106gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(G106gat), .A3(new_n825_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n475_), .A2(G106gat), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n764_), .A2(new_n766_), .A3(new_n794_), .A4(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n822_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n823_), .A2(G106gat), .A3(new_n825_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n825_), .B1(new_n823_), .B2(G106gat), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n822_), .B(new_n831_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n821_), .B1(new_n832_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n831_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT112), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n835_), .A3(new_n820_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(G1339gat));
  NOR2_X1   g640(.A1(new_n663_), .A2(new_n450_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n475_), .A3(new_n661_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846_));
  INV_X1    g645(.A(new_n617_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT12), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n593_), .B2(new_n540_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n587_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n623_), .B(new_n624_), .C1(new_n850_), .C2(new_n580_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT67), .B1(new_n589_), .B2(new_n626_), .ZN(new_n852_));
  OAI22_X1  g651(.A1(new_n847_), .A2(new_n849_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n846_), .B1(new_n853_), .B2(new_n621_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n631_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n628_), .A2(new_n630_), .A3(KEYINPUT55), .A4(new_n620_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n845_), .B(new_n636_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n495_), .B(new_n502_), .C1(new_n498_), .C2(new_n500_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n496_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n510_), .A3(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n512_), .A2(new_n862_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n863_), .A2(new_n639_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n859_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n620_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n631_), .B1(new_n866_), .B2(new_n846_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n638_), .B1(new_n867_), .B2(new_n857_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n845_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n844_), .B1(new_n865_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n636_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT56), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n872_), .A2(KEYINPUT58), .A3(new_n859_), .A4(new_n864_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n727_), .A3(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n871_), .A2(KEYINPUT113), .A3(KEYINPUT56), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n845_), .B1(new_n868_), .B2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n513_), .A2(new_n639_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n875_), .A2(new_n877_), .A3(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n640_), .A2(new_n642_), .A3(new_n863_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n658_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n874_), .B1(new_n882_), .B2(KEYINPUT57), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n884_), .B(new_n658_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n556_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n614_), .B(new_n514_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT54), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n843_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT114), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n887_), .B(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n881_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n871_), .A2(KEYINPUT113), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n878_), .B1(new_n896_), .B2(new_n845_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n897_), .B2(new_n875_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n884_), .B1(new_n898_), .B2(new_n658_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n882_), .A2(KEYINPUT57), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n874_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n894_), .B1(new_n901_), .B2(new_n556_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n892_), .B(KEYINPUT59), .C1(new_n902_), .C2(new_n843_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n886_), .A2(new_n888_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n307_), .A2(new_n399_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT115), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(new_n906_), .A3(new_n842_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n843_), .A2(KEYINPUT115), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n890_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(KEYINPUT116), .B1(new_n904_), .B2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n912_), .B(new_n909_), .C1(new_n886_), .C2(new_n888_), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n891_), .B(new_n903_), .C1(new_n911_), .C2(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G113gat), .B1(new_n914_), .B2(new_n514_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n889_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n514_), .A2(G113gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(G1340gat));
  OR2_X1    g717(.A1(new_n911_), .A2(new_n913_), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n919_), .A2(new_n645_), .A3(new_n903_), .A4(new_n891_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n920_), .A2(KEYINPUT118), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT117), .B(G120gat), .Z(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n923_), .B1(new_n920_), .B2(KEYINPUT118), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n765_), .B2(KEYINPUT60), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(KEYINPUT60), .B2(new_n922_), .ZN(new_n926_));
  OAI22_X1  g725(.A1(new_n921_), .A2(new_n924_), .B1(new_n916_), .B2(new_n926_), .ZN(G1341gat));
  OAI21_X1  g726(.A(G127gat), .B1(new_n914_), .B2(new_n556_), .ZN(new_n928_));
  OR3_X1    g727(.A1(new_n916_), .A2(G127gat), .A3(new_n556_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n928_), .A2(KEYINPUT119), .A3(new_n929_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1342gat));
  INV_X1    g733(.A(G134gat), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n914_), .A2(new_n935_), .A3(new_n719_), .ZN(new_n936_));
  AOI21_X1  g735(.A(G134gat), .B1(new_n889_), .B2(new_n659_), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT120), .Z(new_n938_));
  NOR2_X1   g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1343gat));
  AOI211_X1 g738(.A(new_n475_), .B(new_n423_), .C1(new_n886_), .C2(new_n888_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n399_), .A2(new_n450_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n514_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(new_n206_), .ZN(G1344gat));
  NOR2_X1   g743(.A1(new_n942_), .A2(new_n765_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(new_n207_), .ZN(G1345gat));
  NAND3_X1  g745(.A1(new_n940_), .A2(new_n799_), .A3(new_n941_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(KEYINPUT121), .ZN(new_n948_));
  XNOR2_X1  g747(.A(KEYINPUT61), .B(G155gat), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n948_), .B(new_n949_), .ZN(G1346gat));
  OAI21_X1  g749(.A(G162gat), .B1(new_n942_), .B2(new_n719_), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n680_), .A2(G162gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n942_), .B2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n953_), .B(new_n954_), .ZN(G1347gat));
  INV_X1    g754(.A(G169gat), .ZN(new_n956_));
  NOR4_X1   g755(.A1(new_n902_), .A2(new_n307_), .A3(new_n661_), .A4(new_n451_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n956_), .B1(new_n957_), .B2(new_n513_), .ZN(new_n958_));
  OR2_X1    g757(.A1(new_n958_), .A2(KEYINPUT62), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n957_), .A2(new_n323_), .A3(new_n513_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n958_), .A2(KEYINPUT62), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n959_), .A2(new_n960_), .A3(new_n961_), .ZN(G1348gat));
  XNOR2_X1  g761(.A(KEYINPUT123), .B(G176gat), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n324_), .A2(KEYINPUT123), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n957_), .A2(new_n645_), .ZN(new_n965_));
  MUX2_X1   g764(.A(new_n963_), .B(new_n964_), .S(new_n965_), .Z(G1349gat));
  NAND2_X1  g765(.A1(new_n957_), .A2(new_n799_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n967_), .A2(new_n335_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n968_), .B1(new_n315_), .B2(new_n967_), .ZN(G1350gat));
  NAND2_X1  g768(.A1(new_n659_), .A2(new_n336_), .ZN(new_n970_));
  XOR2_X1   g769(.A(new_n970_), .B(KEYINPUT124), .Z(new_n971_));
  NAND2_X1  g770(.A1(new_n957_), .A2(new_n971_), .ZN(new_n972_));
  AND2_X1   g771(.A1(new_n957_), .A2(new_n727_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n973_), .B2(new_n316_), .ZN(G1351gat));
  NOR2_X1   g773(.A1(new_n661_), .A2(new_n449_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n940_), .A2(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n940_), .A2(KEYINPUT125), .A3(new_n975_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n978_), .A2(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n980_), .A2(new_n513_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g781(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n980_), .A2(new_n645_), .A3(new_n983_), .ZN(new_n984_));
  AND2_X1   g783(.A1(new_n978_), .A2(new_n979_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n985_), .A2(new_n765_), .ZN(new_n986_));
  XOR2_X1   g785(.A(KEYINPUT126), .B(G204gat), .Z(new_n987_));
  OAI21_X1  g786(.A(new_n984_), .B1(new_n986_), .B2(new_n987_), .ZN(G1353gat));
  XNOR2_X1  g787(.A(KEYINPUT63), .B(G211gat), .ZN(new_n989_));
  AOI211_X1 g788(.A(new_n556_), .B(new_n989_), .C1(new_n978_), .C2(new_n979_), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n980_), .A2(new_n799_), .ZN(new_n991_));
  NOR2_X1   g790(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n992_));
  AOI21_X1  g791(.A(new_n990_), .B1(new_n991_), .B2(new_n992_), .ZN(G1354gat));
  AND3_X1   g792(.A1(new_n980_), .A2(G218gat), .A3(new_n727_), .ZN(new_n994_));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995_));
  OAI21_X1  g794(.A(new_n995_), .B1(new_n985_), .B2(new_n680_), .ZN(new_n996_));
  AOI21_X1  g795(.A(new_n680_), .B1(new_n978_), .B2(new_n979_), .ZN(new_n997_));
  AOI21_X1  g796(.A(G218gat), .B1(new_n997_), .B2(KEYINPUT127), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n994_), .B1(new_n996_), .B2(new_n998_), .ZN(G1355gat));
endmodule


