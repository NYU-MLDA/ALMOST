//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G106gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT9), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n208_), .A2(new_n211_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n205_), .A2(new_n207_), .A3(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G85gat), .B(G92gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n213_), .A2(new_n215_), .ZN(new_n223_));
  AOI211_X1 g022(.A(KEYINPUT8), .B(new_n218_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n214_), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n219_), .B(new_n229_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n225_), .B1(new_n232_), .B2(new_n206_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n217_), .B1(new_n224_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(KEYINPUT67), .B(new_n217_), .C1(new_n224_), .C2(new_n233_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G29gat), .B(G36gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G43gat), .B(G50gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT15), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n236_), .A2(new_n237_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n205_), .A2(new_n207_), .A3(new_n216_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n232_), .A2(new_n206_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT8), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n232_), .A2(new_n225_), .A3(new_n206_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n244_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n240_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G232gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n242_), .A2(new_n243_), .A3(new_n249_), .A4(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n242_), .A2(new_n243_), .A3(new_n249_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n252_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT35), .B1(new_n242_), .B2(new_n249_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n254_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G190gat), .B(G218gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT69), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G134gat), .B(G162gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT36), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n242_), .A2(new_n249_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n255_), .B(new_n252_), .C1(new_n266_), .C2(KEYINPUT35), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT36), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n262_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n269_), .A3(new_n254_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n264_), .A2(new_n265_), .A3(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT37), .B1(new_n264_), .B2(new_n265_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n202_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT37), .ZN(new_n274_));
  INV_X1    g073(.A(new_n263_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n267_), .B2(new_n254_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n274_), .B1(new_n276_), .B2(KEYINPUT70), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n264_), .A2(new_n270_), .A3(new_n265_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(KEYINPUT71), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n273_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n270_), .B1(new_n264_), .B2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n276_), .A2(KEYINPUT72), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n274_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G183gat), .B(G211gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT76), .ZN(new_n288_));
  XOR2_X1   g087(.A(G127gat), .B(G155gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT78), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G57gat), .B(G64gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G71gat), .B(G78gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(KEYINPUT11), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(KEYINPUT11), .ZN(new_n299_));
  INV_X1    g098(.A(new_n297_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n296_), .A2(KEYINPUT11), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n298_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(G231gat), .A2(G233gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G8gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT73), .Z(new_n309_));
  XNOR2_X1  g108(.A(G15gat), .B(G22gat), .ZN(new_n310_));
  INV_X1    g109(.A(G1gat), .ZN(new_n311_));
  INV_X1    g110(.A(G8gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT14), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n308_), .B(KEYINPUT73), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n314_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n307_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n307_), .A2(new_n319_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n295_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n307_), .B(new_n319_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n292_), .B(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n286_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT80), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT90), .Z(new_n332_));
  INV_X1    g131(.A(G197gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(G204gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT89), .ZN(new_n335_));
  INV_X1    g134(.A(G204gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n336_), .A2(G197gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n332_), .A2(KEYINPUT21), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n331_), .B(KEYINPUT90), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT21), .B1(new_n337_), .B2(new_n334_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n341_), .B(new_n342_), .C1(new_n339_), .C2(KEYINPUT21), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G169gat), .ZN(new_n346_));
  INV_X1    g145(.A(G183gat), .ZN(new_n347_));
  INV_X1    g146(.A(G190gat), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT23), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(G183gat), .B2(G190gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n346_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n355_));
  INV_X1    g154(.A(G169gat), .ZN(new_n356_));
  INV_X1    g155(.A(G176gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT24), .B1(new_n356_), .B2(new_n357_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT25), .B(G183gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT26), .B1(new_n364_), .B2(new_n348_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT26), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT82), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n363_), .A2(new_n370_), .A3(new_n365_), .A4(new_n367_), .ZN(new_n371_));
  AOI211_X1 g170(.A(KEYINPUT84), .B(new_n362_), .C1(new_n369_), .C2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n351_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT23), .B1(new_n347_), .B2(new_n348_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT85), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n349_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT24), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(new_n360_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n362_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n344_), .B(new_n354_), .C1(new_n372_), .C2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n340_), .A2(new_n343_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n346_), .B(KEYINPUT92), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n374_), .A2(new_n376_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n349_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n353_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT93), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT93), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n377_), .B2(new_n353_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n385_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT26), .B(G190gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n352_), .B1(new_n363_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n360_), .ZN(new_n396_));
  XOR2_X1   g195(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n397_));
  OR2_X1    g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n396_), .B(new_n397_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n395_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n384_), .B1(new_n393_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n383_), .A2(KEYINPUT20), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT19), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n393_), .A2(new_n400_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(new_n344_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n404_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n354_), .B1(new_n382_), .B2(new_n372_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n384_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n408_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n405_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT18), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n405_), .A2(new_n417_), .A3(new_n412_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT3), .ZN(new_n425_));
  INV_X1    g224(.A(G141gat), .ZN(new_n426_));
  INV_X1    g225(.A(G148gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G141gat), .A2(G148gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT2), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n428_), .A2(new_n431_), .A3(new_n432_), .A4(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(G155gat), .A2(G162gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G155gat), .A2(G162gat), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G141gat), .B(G148gat), .Z(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(KEYINPUT1), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n435_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n436_), .A2(KEYINPUT1), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n439_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n438_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT95), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G127gat), .B(G134gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G113gat), .B(G120gat), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n448_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n446_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n438_), .A2(new_n443_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(KEYINPUT95), .ZN(new_n454_));
  INV_X1    g253(.A(new_n451_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT4), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n444_), .A2(KEYINPUT4), .A3(new_n451_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n424_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n446_), .A2(new_n451_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n454_), .A2(new_n455_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n424_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G29gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G85gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT0), .B(G57gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n466_), .B(new_n467_), .Z(new_n468_));
  NOR3_X1   g267(.A1(new_n460_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n424_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT4), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n473_), .B2(new_n458_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n470_), .B1(new_n474_), .B2(new_n463_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n469_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n402_), .A2(new_n404_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n409_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n417_), .B(KEYINPUT97), .ZN(new_n480_));
  OAI211_X1 g279(.A(KEYINPUT27), .B(new_n420_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n423_), .A2(new_n476_), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n344_), .B1(KEYINPUT29), .B2(new_n453_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n453_), .A2(KEYINPUT29), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n484_), .B(KEYINPUT28), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n483_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G228gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(G78gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(new_n228_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G22gat), .B(G50gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n486_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n451_), .B(KEYINPUT31), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n410_), .A2(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(KEYINPUT30), .B(new_n354_), .C1(new_n382_), .C2(new_n372_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G71gat), .B(G99gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT87), .ZN(new_n500_));
  INV_X1    g299(.A(G15gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G227gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n497_), .A2(new_n498_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT86), .B(G43gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n504_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n380_), .A2(new_n381_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n372_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n379_), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT30), .B1(new_n513_), .B2(new_n354_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n498_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n510_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n497_), .A2(new_n504_), .A3(new_n498_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n507_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT88), .B1(new_n509_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n508_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n516_), .A2(new_n507_), .A3(new_n517_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n495_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n495_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n493_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n522_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n494_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n493_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n525_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n482_), .B1(new_n527_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT96), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n405_), .A2(new_n535_), .A3(new_n412_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n417_), .A2(KEYINPUT32), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n479_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n413_), .B2(new_n535_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n476_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n468_), .B1(new_n460_), .B2(new_n464_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT33), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n457_), .A2(new_n424_), .A3(new_n459_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n452_), .A2(new_n456_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n545_), .B(new_n470_), .C1(new_n424_), .C2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n475_), .A2(KEYINPUT33), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n421_), .B2(KEYINPUT94), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n419_), .A2(new_n551_), .A3(new_n420_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n541_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n530_), .A2(new_n493_), .A3(new_n525_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n534_), .A2(new_n556_), .ZN(new_n557_));
  OAI211_X1 g356(.A(KEYINPUT12), .B(new_n298_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n236_), .A2(new_n237_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n303_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n234_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n248_), .B2(new_n303_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n303_), .B(new_n217_), .C1(new_n224_), .C2(new_n233_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT65), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n246_), .A2(new_n247_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT65), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n571_), .A2(new_n572_), .A3(new_n217_), .A4(new_n303_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n573_), .A3(new_n562_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n565_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT66), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n574_), .A2(KEYINPUT66), .A3(new_n565_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n568_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G120gat), .B(G148gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G176gat), .B(G204gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n581_), .B(new_n582_), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n584_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(KEYINPUT13), .A3(new_n586_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n241_), .A2(new_n319_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n316_), .A2(new_n318_), .A3(new_n240_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n594_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n316_), .A2(new_n318_), .A3(new_n240_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n240_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(G113gat), .B(G141gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n595_), .A2(new_n599_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n591_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n330_), .A2(new_n557_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n476_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n609_), .A2(new_n311_), .A3(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(KEYINPUT38), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n607_), .A2(KEYINPUT98), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n591_), .A2(new_n616_), .A3(new_n606_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n284_), .B1(new_n534_), .B2(new_n556_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(new_n328_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n311_), .B1(new_n622_), .B2(new_n610_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n611_), .B2(KEYINPUT38), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n614_), .A2(new_n624_), .ZN(G1324gat));
  NAND2_X1  g424(.A1(new_n423_), .A2(new_n481_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n609_), .A2(new_n312_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n621_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n312_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT100), .B1(new_n621_), .B2(new_n628_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n627_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT40), .B(new_n627_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1325gat));
  NOR2_X1   g439(.A1(new_n524_), .A2(new_n526_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n609_), .A2(new_n501_), .A3(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT101), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n501_), .B1(new_n622_), .B2(new_n642_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT41), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT41), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n647_), .A3(new_n648_), .ZN(G1326gat));
  OAI21_X1  g448(.A(G22gat), .B1(new_n621_), .B2(new_n493_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT42), .ZN(new_n651_));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n609_), .A2(new_n652_), .A3(new_n531_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1327gat));
  NOR2_X1   g453(.A1(new_n618_), .A2(new_n328_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n273_), .A2(new_n279_), .B1(new_n274_), .B2(new_n284_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n656_), .B1(new_n533_), .B2(new_n555_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(KEYINPUT102), .A3(KEYINPUT43), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT43), .B1(new_n657_), .B2(KEYINPUT102), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT44), .B(new_n655_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n610_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G29gat), .ZN(new_n666_));
  INV_X1    g465(.A(new_n284_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n328_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n608_), .B(new_n668_), .C1(new_n533_), .C2(new_n555_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n476_), .A2(G29gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT103), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n669_), .B2(new_n671_), .ZN(G1328gat));
  NAND3_X1  g471(.A1(new_n662_), .A2(new_n626_), .A3(new_n663_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G36gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n669_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n628_), .A2(G36gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n677_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT104), .B1(new_n669_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT45), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n674_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT46), .B1(new_n683_), .B2(KEYINPUT105), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  AOI211_X1 g485(.A(new_n685_), .B(new_n686_), .C1(new_n674_), .C2(new_n682_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n684_), .A2(new_n687_), .ZN(G1329gat));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n689_));
  INV_X1    g488(.A(G43gat), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n641_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n664_), .A2(new_n689_), .A3(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n669_), .A2(new_n641_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(G43gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n662_), .A2(new_n663_), .A3(new_n691_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(KEYINPUT106), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n692_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1330gat));
  AOI21_X1  g499(.A(G50gat), .B1(new_n675_), .B2(new_n531_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n531_), .A2(G50gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n664_), .B2(new_n702_), .ZN(G1331gat));
  NOR2_X1   g502(.A1(new_n591_), .A2(new_n606_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n330_), .A2(new_n557_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(G57gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n610_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n591_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n327_), .A2(new_n606_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n620_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n476_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(G1332gat));
  OAI21_X1  g511(.A(G64gat), .B1(new_n710_), .B2(new_n628_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT48), .ZN(new_n714_));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n705_), .A2(new_n715_), .A3(new_n626_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n710_), .B2(new_n641_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n705_), .A2(new_n721_), .A3(new_n642_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1334gat));
  OAI21_X1  g522(.A(G78gat), .B1(new_n710_), .B2(new_n493_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT50), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n705_), .A2(new_n488_), .A3(new_n531_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1335gat));
  NOR3_X1   g526(.A1(new_n591_), .A2(new_n328_), .A3(new_n606_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n728_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n476_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n668_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n534_), .B2(new_n556_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n704_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n209_), .A3(new_n610_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n730_), .A2(new_n735_), .ZN(G1336gat));
  OAI21_X1  g535(.A(G92gat), .B1(new_n729_), .B2(new_n628_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n210_), .A3(new_n626_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1337gat));
  AND4_X1   g538(.A1(new_n203_), .A2(new_n732_), .A3(new_n642_), .A4(new_n704_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT110), .Z(new_n741_));
  OAI211_X1 g540(.A(new_n642_), .B(new_n728_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT109), .B1(new_n742_), .B2(G99gat), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(KEYINPUT109), .A3(G99gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n741_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(G1338gat));
  NAND3_X1  g546(.A1(new_n734_), .A2(new_n204_), .A3(new_n531_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n749_));
  OAI21_X1  g548(.A(G106gat), .B1(new_n729_), .B2(new_n493_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT52), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT52), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n748_), .B(new_n749_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n750_), .B(KEYINPUT52), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n749_), .B1(new_n755_), .B2(new_n748_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1339gat));
  NAND3_X1  g556(.A1(new_n709_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n286_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n760_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n656_), .B2(new_n758_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n605_), .B1(new_n579_), .B2(new_n584_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n560_), .A2(new_n564_), .A3(new_n570_), .A4(new_n573_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n565_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n560_), .A2(new_n564_), .A3(new_n566_), .A4(KEYINPUT55), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n567_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n769_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT114), .B1(new_n772_), .B2(new_n583_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n766_), .B1(new_n773_), .B2(KEYINPUT56), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n565_), .A2(new_n767_), .B1(new_n567_), .B2(new_n770_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n584_), .B1(new_n775_), .B2(new_n769_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n776_), .A2(KEYINPUT114), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n765_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n776_), .B2(KEYINPUT114), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n773_), .A2(KEYINPUT56), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(KEYINPUT115), .A4(new_n766_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n592_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n597_), .A2(new_n598_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n602_), .B1(new_n784_), .B2(new_n594_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n603_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n587_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n779_), .A2(new_n782_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n667_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n284_), .A2(new_n790_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n788_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n772_), .A2(new_n583_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n586_), .B(new_n786_), .C1(new_n794_), .C2(KEYINPUT56), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n776_), .A2(new_n777_), .ZN(new_n797_));
  OR3_X1    g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n280_), .A2(new_n285_), .A3(new_n798_), .A4(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n791_), .A2(new_n793_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n764_), .B1(new_n801_), .B2(new_n327_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n527_), .A2(new_n476_), .A3(new_n626_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT59), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n800_), .A2(new_n793_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT57), .B1(new_n788_), .B2(new_n667_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n327_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT116), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n327_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n764_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n804_), .A2(KEYINPUT59), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n805_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT117), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n805_), .B(new_n816_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  INV_X1    g616(.A(G113gat), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n605_), .A2(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT118), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n815_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n764_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n808_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n803_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n818_), .B1(new_n824_), .B2(new_n605_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n821_), .A2(new_n825_), .ZN(G1340gat));
  OR2_X1    g625(.A1(new_n814_), .A2(new_n591_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G120gat), .ZN(new_n828_));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n591_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(KEYINPUT60), .B2(new_n829_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n828_), .B1(new_n824_), .B2(new_n831_), .ZN(G1341gat));
  NAND3_X1  g631(.A1(new_n815_), .A2(new_n328_), .A3(new_n817_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G127gat), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n327_), .A2(G127gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n824_), .B2(new_n835_), .ZN(G1342gat));
  XNOR2_X1  g635(.A(KEYINPUT119), .B(G134gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n656_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n815_), .A2(new_n817_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(G134gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n824_), .B2(new_n667_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT120), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n840_), .A2(new_n845_), .A3(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1343gat));
  NOR2_X1   g646(.A1(new_n802_), .A2(new_n532_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n626_), .A2(new_n476_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n605_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(new_n426_), .ZN(G1344gat));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n591_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n427_), .ZN(G1345gat));
  NAND3_X1  g653(.A1(new_n848_), .A2(new_n328_), .A3(new_n849_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT121), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n856_), .B(new_n858_), .ZN(G1346gat));
  NOR2_X1   g658(.A1(new_n850_), .A2(new_n667_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n656_), .A2(G162gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT122), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n860_), .A2(G162gat), .B1(new_n850_), .B2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT123), .ZN(G1347gat));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n628_), .A2(new_n610_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n642_), .A3(new_n493_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n812_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n606_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n865_), .B1(new_n869_), .B2(G169gat), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n869_), .A2(new_n865_), .A3(G169gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(KEYINPUT62), .A3(new_n872_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT22), .B(G169gat), .Z(new_n874_));
  NOR2_X1   g673(.A1(new_n869_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n870_), .B2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n877_), .ZN(G1348gat));
  AOI21_X1  g677(.A(G176gat), .B1(new_n868_), .B2(new_n708_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n867_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n591_), .A2(new_n357_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n823_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT125), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n879_), .A2(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT126), .ZN(G1349gat));
  NOR2_X1   g684(.A1(new_n327_), .A2(new_n363_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n823_), .A2(new_n328_), .A3(new_n880_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n868_), .A2(new_n886_), .B1(new_n347_), .B2(new_n887_), .ZN(G1350gat));
  NAND3_X1  g687(.A1(new_n868_), .A2(new_n284_), .A3(new_n394_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n812_), .A2(new_n286_), .A3(new_n867_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n348_), .ZN(G1351gat));
  NAND2_X1  g690(.A1(new_n848_), .A2(new_n866_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n605_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n333_), .ZN(G1352gat));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n591_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n336_), .ZN(G1353gat));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  AND2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n892_), .A2(new_n327_), .A3(new_n897_), .A4(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n848_), .A2(new_n328_), .A3(new_n866_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n897_), .ZN(G1354gat));
  OAI21_X1  g700(.A(G218gat), .B1(new_n892_), .B2(new_n286_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n667_), .A2(G218gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n892_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT127), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1355gat));
endmodule


