//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n829_, new_n831_, new_n832_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n854_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT83), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(new_n203_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT83), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT84), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT31), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G227gat), .A2(G233gat), .ZN(new_n213_));
  INV_X1    g012(.A(G15gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT30), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT79), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n218_), .B(new_n220_), .C1(new_n226_), .C2(KEYINPUT24), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT24), .B1(new_n224_), .B2(new_n225_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n219_), .B(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT80), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n232_), .A4(new_n225_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT25), .B(G183gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT78), .ZN(new_n235_));
  INV_X1    g034(.A(G190gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n235_), .B1(new_n236_), .B2(KEYINPUT26), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT26), .B(G190gat), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n234_), .B(new_n237_), .C1(new_n238_), .C2(new_n235_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n227_), .A2(new_n231_), .A3(new_n233_), .A4(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n220_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT22), .B(G169gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT82), .B(G176gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n222_), .B2(KEYINPUT22), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n242_), .B(new_n232_), .C1(new_n245_), .C2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G71gat), .B(G99gat), .ZN(new_n250_));
  INV_X1    g049(.A(G43gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n240_), .A2(new_n249_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n240_), .B2(new_n249_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n217_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n240_), .A2(new_n249_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n252_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(new_n216_), .A3(new_n254_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT85), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n212_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n260_), .A3(KEYINPUT85), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT86), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT86), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n257_), .A2(new_n260_), .A3(KEYINPUT85), .A4(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n267_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n257_), .A2(new_n260_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n270_), .A2(KEYINPUT85), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n269_), .B1(new_n271_), .B2(new_n212_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G78gat), .B(G106gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT90), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G211gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(G218gat), .ZN(new_n277_));
  INV_X1    g076(.A(G218gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(G211gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT89), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G197gat), .A2(G204gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G197gat), .A2(G204gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(KEYINPUT21), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  INV_X1    g084(.A(new_n283_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(new_n286_), .B2(new_n281_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n278_), .A2(G211gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n276_), .A2(G218gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT89), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n280_), .A2(new_n284_), .A3(new_n287_), .A4(new_n291_), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n286_), .A2(new_n281_), .A3(new_n285_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n290_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT2), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n301_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT88), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n302_), .A2(new_n305_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n300_), .A2(KEYINPUT1), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n300_), .B1(new_n298_), .B2(KEYINPUT1), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(KEYINPUT87), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT87), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n314_), .B(new_n300_), .C1(new_n298_), .C2(KEYINPUT1), .ZN(new_n315_));
  AOI211_X1 g114(.A(new_n309_), .B(new_n310_), .C1(new_n313_), .C2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(KEYINPUT87), .ZN(new_n317_));
  INV_X1    g116(.A(new_n311_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n310_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT88), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n308_), .B1(new_n316_), .B2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n297_), .B1(new_n322_), .B2(KEYINPUT29), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n324_), .ZN(new_n326_));
  AOI211_X1 g125(.A(new_n297_), .B(new_n326_), .C1(new_n322_), .C2(KEYINPUT29), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n275_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT91), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n319_), .A2(new_n320_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n309_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n319_), .A2(KEYINPUT88), .A3(new_n320_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n307_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G22gat), .B(G50gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT28), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n336_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n297_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n326_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n323_), .A2(new_n324_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(new_n274_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n330_), .A2(new_n339_), .B1(new_n344_), .B2(new_n328_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n328_), .A2(new_n344_), .A3(KEYINPUT91), .A4(new_n339_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n268_), .B(new_n272_), .C1(new_n345_), .C2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n274_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n339_), .B1(new_n349_), .B2(KEYINPUT91), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n328_), .A2(new_n344_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n268_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n263_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n346_), .B(new_n352_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n348_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n210_), .A2(new_n322_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n207_), .A2(new_n204_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n334_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n358_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(KEYINPUT4), .B1(new_n210_), .B2(new_n322_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n361_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(KEYINPUT4), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n365_), .B2(new_n358_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G1gat), .B(G29gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(G57gat), .B(G85gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n366_), .A2(new_n372_), .ZN(new_n373_));
  AOI211_X1 g172(.A(new_n357_), .B(new_n363_), .C1(new_n364_), .C2(KEYINPUT4), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n371_), .B1(new_n374_), .B2(new_n362_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n356_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT98), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n258_), .A2(new_n340_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n243_), .A2(new_n246_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n232_), .B(KEYINPUT93), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT94), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n382_), .A3(KEYINPUT94), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n242_), .A3(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n228_), .A2(new_n230_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n238_), .A2(new_n234_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n233_), .A3(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(new_n297_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT19), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n380_), .A2(KEYINPUT20), .A3(new_n391_), .A4(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT96), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n240_), .A2(new_n297_), .A3(new_n249_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT92), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n397_), .A2(new_n398_), .A3(KEYINPUT20), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n397_), .B2(KEYINPUT20), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n297_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT95), .B1(new_n402_), .B2(new_n394_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n400_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n397_), .A2(new_n398_), .A3(KEYINPUT20), .ZN(new_n405_));
  INV_X1    g204(.A(new_n401_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT95), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n393_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n396_), .B1(new_n403_), .B2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G8gat), .B(G36gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT18), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G64gat), .B(G92gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  OAI21_X1  g213(.A(new_n379_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n395_), .B(KEYINPUT96), .Z(new_n416_));
  NOR3_X1   g215(.A1(new_n402_), .A2(KEYINPUT95), .A3(new_n394_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n408_), .B1(new_n407_), .B2(new_n393_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n414_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(KEYINPUT98), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n415_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT27), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n410_), .A2(new_n414_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT97), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n410_), .A2(KEYINPUT97), .A3(new_n414_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n422_), .A2(new_n423_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n380_), .A2(KEYINPUT20), .A3(new_n391_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n393_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n407_), .B2(new_n393_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n420_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n432_), .A2(KEYINPUT101), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(KEYINPUT101), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n424_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT27), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n378_), .B1(new_n428_), .B2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n345_), .A2(new_n347_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n353_), .A2(new_n354_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT33), .B1(new_n366_), .B2(new_n372_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n442_), .B(new_n371_), .C1(new_n374_), .C2(new_n362_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n365_), .A2(new_n358_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n372_), .B1(new_n364_), .B2(new_n357_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT100), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n445_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT100), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n447_), .B(new_n448_), .C1(new_n358_), .C2(new_n365_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n441_), .A2(new_n443_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n422_), .A2(new_n426_), .A3(new_n427_), .A4(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n414_), .A2(KEYINPUT32), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n431_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n376_), .B(new_n453_), .C1(new_n419_), .C2(new_n452_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n440_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n437_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G57gat), .B(G64gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT11), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT65), .ZN(new_n459_));
  XOR2_X1   g258(.A(G71gat), .B(G78gat), .Z(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(KEYINPUT11), .B2(new_n457_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n459_), .B(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT10), .B(G99gat), .Z(new_n463_));
  INV_X1    g262(.A(G106gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G85gat), .B(G92gat), .Z(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT9), .ZN(new_n467_));
  INV_X1    g266(.A(G85gat), .ZN(new_n468_));
  INV_X1    g267(.A(G92gat), .ZN(new_n469_));
  OR3_X1    g268(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT9), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT6), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(G99gat), .A3(G106gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n465_), .A2(new_n467_), .A3(new_n470_), .A4(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT64), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n473_), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n471_), .A2(KEYINPUT6), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n472_), .A2(new_n474_), .A3(KEYINPUT64), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n481_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n477_), .B1(new_n487_), .B2(new_n466_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n466_), .A2(new_n477_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n475_), .B2(new_n486_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n476_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n462_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n462_), .A2(new_n491_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT12), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G230gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(KEYINPUT66), .B(new_n476_), .C1(new_n488_), .C2(new_n490_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n498_), .A2(KEYINPUT12), .A3(new_n462_), .A4(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n496_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n492_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n502_), .B1(new_n503_), .B2(new_n493_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G176gat), .B(G204gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT68), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G120gat), .B(G148gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n505_), .B(new_n511_), .Z(new_n512_));
  INV_X1    g311(.A(KEYINPUT13), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n513_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517_));
  INV_X1    g316(.A(G1gat), .ZN(new_n518_));
  INV_X1    g317(.A(G8gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G1gat), .B(G8gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G29gat), .B(G36gat), .Z(new_n526_));
  XOR2_X1   g325(.A(G43gat), .B(G50gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT15), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(KEYINPUT75), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n528_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n525_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(KEYINPUT75), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n531_), .A2(new_n532_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n525_), .B(new_n533_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n532_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G113gat), .B(G141gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT76), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G169gat), .B(G197gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  NAND3_X1  g342(.A1(new_n536_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT77), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT77), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n536_), .A2(new_n539_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n543_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n545_), .A2(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n516_), .A2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n456_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G134gat), .B(G162gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n498_), .A2(new_n529_), .A3(new_n499_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT34), .Z(new_n558_));
  INV_X1    g357(.A(KEYINPUT35), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n528_), .B(new_n476_), .C1(new_n488_), .C2(new_n490_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n559_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT70), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n556_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n565_), .B1(new_n556_), .B2(KEYINPUT69), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT69), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n498_), .A2(new_n570_), .A3(new_n529_), .A4(new_n499_), .ZN(new_n571_));
  AOI211_X1 g370(.A(new_n568_), .B(new_n561_), .C1(new_n569_), .C2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n556_), .A2(KEYINPUT69), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n571_), .A3(new_n566_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT71), .B1(new_n574_), .B2(new_n560_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n555_), .B(new_n567_), .C1(new_n572_), .C2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(KEYINPUT72), .B(new_n567_), .C1(new_n572_), .C2(new_n575_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n555_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n552_), .A2(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n577_), .A2(new_n552_), .A3(new_n578_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT37), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(new_n552_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n578_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n577_), .A2(new_n552_), .A3(new_n578_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n581_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n525_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(new_n462_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT16), .ZN(new_n594_));
  XOR2_X1   g393(.A(G183gat), .B(G211gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n597_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n592_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n599_), .B2(new_n592_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n589_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n551_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n518_), .A3(new_n376_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT38), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n579_), .A2(new_n580_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n602_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n551_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G1gat), .B1(new_n612_), .B2(new_n377_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n613_), .ZN(G1324gat));
  NAND2_X1  g413(.A1(new_n428_), .A2(new_n436_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G8gat), .B1(new_n612_), .B2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT39), .ZN(new_n617_));
  INV_X1    g416(.A(new_n615_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n606_), .A2(new_n519_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g420(.A(new_n439_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n606_), .A2(new_n214_), .A3(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT102), .Z(new_n624_));
  OAI21_X1  g423(.A(G15gat), .B1(new_n612_), .B2(new_n439_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT41), .Z(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(G1326gat));
  OAI21_X1  g426(.A(G22gat), .B1(new_n612_), .B2(new_n438_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT42), .ZN(new_n629_));
  INV_X1    g428(.A(G22gat), .ZN(new_n630_));
  INV_X1    g429(.A(new_n438_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n606_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(G1327gat));
  NOR2_X1   g432(.A1(new_n609_), .A2(new_n603_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n551_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n376_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n588_), .B2(KEYINPUT103), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n588_), .B1(new_n437_), .B2(new_n455_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI221_X1 g441(.A(new_n588_), .B1(KEYINPUT103), .B2(new_n639_), .C1(new_n437_), .C2(new_n455_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n550_), .A2(new_n602_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT44), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n648_), .B(new_n645_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n637_), .B1(new_n650_), .B2(new_n376_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n638_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  NAND2_X1  g454(.A1(new_n644_), .A2(new_n646_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n648_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n646_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n618_), .A4(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G36gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n658_), .B1(new_n650_), .B2(new_n618_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT106), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n657_), .A2(new_n618_), .A3(new_n659_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT105), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(G36gat), .A4(new_n660_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n615_), .A2(G36gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n636_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT107), .B1(new_n635_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT45), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n668_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n668_), .A2(KEYINPUT46), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1329gat));
  AOI21_X1  g479(.A(G43gat), .B1(new_n636_), .B2(new_n622_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n439_), .A2(new_n251_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n650_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(G1330gat));
  AOI21_X1  g484(.A(G50gat), .B1(new_n636_), .B2(new_n631_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n631_), .A2(G50gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n650_), .B2(new_n687_), .ZN(G1331gat));
  INV_X1    g487(.A(new_n516_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n549_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n456_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n611_), .ZN(new_n693_));
  INV_X1    g492(.A(G57gat), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n377_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n605_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n377_), .B1(new_n696_), .B2(KEYINPUT109), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n697_), .B1(KEYINPUT109), .B2(new_n696_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n695_), .B1(new_n698_), .B2(new_n694_), .ZN(G1332gat));
  OAI21_X1  g498(.A(G64gat), .B1(new_n693_), .B2(new_n615_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT48), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n615_), .A2(G64gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n696_), .B2(new_n702_), .ZN(G1333gat));
  NAND3_X1  g502(.A1(new_n692_), .A2(new_n622_), .A3(new_n611_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT49), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(G71gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n704_), .B2(G71gat), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n439_), .A2(G71gat), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT110), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n707_), .A2(new_n708_), .B1(new_n696_), .B2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT111), .Z(G1334gat));
  OAI21_X1  g511(.A(G78gat), .B1(new_n693_), .B2(new_n438_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT50), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n438_), .A2(G78gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n696_), .B2(new_n715_), .ZN(G1335gat));
  NAND3_X1  g515(.A1(new_n644_), .A2(new_n602_), .A3(new_n691_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G85gat), .B1(new_n717_), .B2(new_n377_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n692_), .A2(new_n634_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n468_), .A3(new_n376_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1336gat));
  OAI21_X1  g521(.A(G92gat), .B1(new_n717_), .B2(new_n615_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n469_), .A3(new_n618_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1337gat));
  NAND2_X1  g524(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n622_), .A2(new_n463_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n719_), .B2(new_n727_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n717_), .A2(new_n439_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G99gat), .ZN(new_n730_));
  NOR2_X1   g529(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(G1338gat));
  NOR2_X1   g531(.A1(new_n717_), .A2(new_n438_), .ZN(new_n733_));
  OR3_X1    g532(.A1(new_n733_), .A2(KEYINPUT113), .A3(new_n464_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT113), .B1(new_n733_), .B2(new_n464_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(KEYINPUT52), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT113), .B(new_n737_), .C1(new_n733_), .C2(new_n464_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n720_), .A2(new_n464_), .A3(new_n631_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g540(.A1(new_n618_), .A2(new_n377_), .A3(new_n355_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n545_), .A2(new_n546_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n505_), .A2(new_n511_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n543_), .B1(new_n537_), .B2(new_n532_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n747_), .A2(KEYINPUT115), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n531_), .A2(new_n538_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(KEYINPUT115), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n744_), .A2(new_n746_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n501_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n495_), .A2(new_n500_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n502_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT114), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n755_), .A2(new_n758_), .A3(new_n502_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n501_), .A2(new_n753_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n754_), .A2(new_n757_), .A3(new_n759_), .A4(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n511_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT56), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(KEYINPUT56), .A3(new_n511_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n752_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT58), .B1(new_n766_), .B2(KEYINPUT116), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n764_), .A2(new_n765_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n768_), .B(new_n769_), .C1(new_n770_), .C2(new_n752_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n767_), .A2(new_n771_), .A3(new_n588_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n764_), .A2(new_n765_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n549_), .A2(new_n745_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n744_), .A2(new_n751_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(new_n512_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT57), .B(new_n609_), .C1(new_n775_), .C2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n777_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(new_n610_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n772_), .A2(new_n778_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n602_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n516_), .A2(new_n690_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n589_), .A2(new_n784_), .A3(new_n603_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT54), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n589_), .A2(new_n784_), .A3(new_n787_), .A4(new_n603_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n743_), .B1(new_n783_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(G113gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n690_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n742_), .A2(new_n793_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(KEYINPUT119), .B2(new_n743_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n782_), .A2(new_n602_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT59), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT117), .B1(new_n790_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(KEYINPUT59), .C1(new_n798_), .C2(new_n743_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n799_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT120), .B(new_n799_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n549_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n792_), .B1(new_n808_), .B2(new_n791_), .ZN(G1340gat));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n689_), .B2(KEYINPUT60), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n790_), .B(new_n811_), .C1(KEYINPUT60), .C2(new_n810_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n804_), .A2(new_n516_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n810_), .ZN(G1341gat));
  AOI21_X1  g613(.A(G127gat), .B1(new_n790_), .B2(new_n603_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n806_), .A2(new_n807_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n603_), .A2(G127gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT121), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n815_), .B1(new_n816_), .B2(new_n818_), .ZN(G1342gat));
  AOI21_X1  g618(.A(G134gat), .B1(new_n790_), .B2(new_n610_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT122), .Z(new_n821_));
  AND2_X1   g620(.A1(new_n588_), .A2(G134gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n816_), .B2(new_n822_), .ZN(G1343gat));
  NOR2_X1   g622(.A1(new_n798_), .A2(new_n348_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n376_), .A3(new_n615_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n549_), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g626(.A1(new_n825_), .A2(new_n689_), .ZN(new_n828_));
  XOR2_X1   g627(.A(KEYINPUT123), .B(G148gat), .Z(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1345gat));
  NOR2_X1   g629(.A1(new_n825_), .A2(new_n602_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT61), .B(G155gat), .Z(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1346gat));
  OAI21_X1  g632(.A(G162gat), .B1(new_n825_), .B2(new_n589_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n609_), .A2(G162gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n825_), .B2(new_n835_), .ZN(G1347gat));
  NOR2_X1   g635(.A1(new_n798_), .A2(new_n631_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n615_), .A2(new_n376_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n622_), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT124), .Z(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n690_), .A3(new_n243_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n840_), .A2(new_n690_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT125), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n837_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n844_), .B1(new_n847_), .B2(G169gat), .ZN(new_n848_));
  AOI211_X1 g647(.A(KEYINPUT62), .B(new_n222_), .C1(new_n846_), .C2(new_n837_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n843_), .B1(new_n848_), .B2(new_n849_), .ZN(G1348gat));
  NAND2_X1  g649(.A1(new_n842_), .A2(new_n516_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n223_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n246_), .B2(new_n851_), .ZN(G1349gat));
  NOR2_X1   g652(.A1(new_n841_), .A2(new_n602_), .ZN(new_n854_));
  MUX2_X1   g653(.A(G183gat), .B(new_n234_), .S(new_n854_), .Z(G1350gat));
  OAI21_X1  g654(.A(G190gat), .B1(new_n841_), .B2(new_n589_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n610_), .A2(new_n238_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n841_), .B2(new_n857_), .ZN(G1351gat));
  NAND2_X1  g657(.A1(new_n824_), .A2(new_n838_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n549_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n689_), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(G204gat), .Z(G1353gat));
  NOR2_X1   g662(.A1(new_n859_), .A2(new_n602_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n864_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT63), .B(G211gat), .Z(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n864_), .B2(new_n866_), .ZN(G1354gat));
  XOR2_X1   g666(.A(KEYINPUT126), .B(G218gat), .Z(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n859_), .B2(new_n609_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n589_), .A2(new_n868_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n859_), .B2(new_n870_), .ZN(new_n871_));
  XOR2_X1   g670(.A(new_n871_), .B(KEYINPUT127), .Z(G1355gat));
endmodule


