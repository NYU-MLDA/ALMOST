//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT19), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT23), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT76), .B(KEYINPUT23), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(new_n210_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT22), .B(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT95), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT95), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n218_), .A2(new_n222_), .A3(new_n219_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n215_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT92), .ZN(new_n226_));
  INV_X1    g025(.A(G169gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n217_), .A3(KEYINPUT75), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n229_), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT92), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n219_), .A2(new_n231_), .A3(KEYINPUT24), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n226_), .A2(new_n228_), .A3(new_n230_), .A4(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT25), .B(G183gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT26), .B(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n233_), .A2(KEYINPUT93), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n210_), .ZN(new_n238_));
  AND2_X1   g037(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n239_));
  NOR2_X1   g038(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT24), .B1(new_n228_), .B2(new_n230_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT94), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n242_), .B1(new_n212_), .B2(new_n238_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n228_), .A2(new_n230_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT24), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT94), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n237_), .A2(new_n246_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT93), .B1(new_n233_), .B2(new_n236_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n224_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G197gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT85), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G197gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n259_), .A3(G204gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT87), .B1(new_n256_), .B2(G204gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT87), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n257_), .A2(new_n259_), .A3(new_n264_), .A4(G204gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n263_), .A2(KEYINPUT21), .A3(new_n265_), .A4(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT21), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT85), .B(G197gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n261_), .B1(new_n270_), .B2(G204gat), .ZN(new_n271_));
  AND4_X1   g070(.A1(new_n264_), .A2(new_n257_), .A3(new_n259_), .A4(G204gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n269_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n266_), .ZN(new_n274_));
  INV_X1    g073(.A(G204gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n257_), .A2(new_n259_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n269_), .B1(G197gat), .B2(G204gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(KEYINPUT86), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT86), .B1(new_n276_), .B2(new_n277_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n268_), .B1(new_n274_), .B2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT20), .B1(new_n255_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT100), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n236_), .B1(new_n248_), .B2(new_n225_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n285_), .A2(new_n213_), .A3(new_n245_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(G176gat), .B1(new_n227_), .B2(KEYINPUT22), .ZN(new_n288_));
  OR2_X1    g087(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n289_));
  NAND2_X1  g088(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n227_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n288_), .B1(new_n291_), .B2(KEYINPUT78), .ZN(new_n292_));
  AND2_X1   g091(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n293_));
  NOR2_X1   g092(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n294_));
  OAI211_X1 g093(.A(KEYINPUT78), .B(G169gat), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(KEYINPUT79), .B(new_n219_), .C1(new_n292_), .C2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n244_), .A2(new_n214_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n219_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n288_), .ZN(new_n302_));
  OAI21_X1  g101(.A(G169gat), .B1(new_n293_), .B2(new_n294_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n301_), .B1(new_n305_), .B2(new_n295_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(KEYINPUT79), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n287_), .B1(new_n300_), .B2(new_n307_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n283_), .A2(new_n284_), .B1(new_n308_), .B2(new_n282_), .ZN(new_n309_));
  AND4_X1   g108(.A1(KEYINPUT21), .A2(new_n263_), .A3(new_n265_), .A4(new_n267_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n263_), .A2(new_n265_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n267_), .B1(new_n311_), .B2(new_n269_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n280_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n278_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n310_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n315_), .B(new_n224_), .C1(new_n254_), .C2(new_n253_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(KEYINPUT100), .A3(KEYINPUT20), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n209_), .B1(new_n309_), .B2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n315_), .B(new_n287_), .C1(new_n307_), .C2(new_n300_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n255_), .A2(new_n282_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(KEYINPUT20), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n208_), .B(KEYINPUT91), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n206_), .B1(new_n318_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(new_n322_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n308_), .A2(new_n282_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n326_), .A2(KEYINPUT20), .A3(new_n209_), .A4(new_n316_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n205_), .A3(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(KEYINPUT27), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n298_), .B1(new_n306_), .B2(KEYINPUT79), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n219_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n286_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n209_), .B1(new_n334_), .B2(new_n315_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(new_n283_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n322_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT20), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n255_), .B2(new_n282_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n339_), .B2(new_n319_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n206_), .B1(new_n336_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n328_), .A3(KEYINPUT96), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT27), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT96), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n344_), .B(new_n206_), .C1(new_n336_), .C2(new_n340_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n329_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G113gat), .B(G120gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT82), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT82), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n349_), .A2(new_n350_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n349_), .A2(new_n350_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G141gat), .B(G148gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(KEYINPUT1), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n360_));
  INV_X1    g159(.A(new_n357_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n359_), .A2(KEYINPUT83), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n363_), .B(new_n357_), .C1(new_n358_), .C2(KEYINPUT1), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n356_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366_));
  INV_X1    g165(.A(G141gat), .ZN(new_n367_));
  INV_X1    g166(.A(G148gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .A4(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n358_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n374_), .A2(new_n357_), .A3(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n351_), .B(new_n355_), .C1(new_n365_), .C2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n357_), .A3(new_n375_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n349_), .B(new_n350_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n359_), .A2(KEYINPUT83), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n361_), .A2(new_n360_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n380_), .A2(new_n364_), .A3(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n378_), .B(new_n379_), .C1(new_n382_), .C2(new_n356_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n377_), .A2(KEYINPUT4), .A3(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n378_), .B1(new_n382_), .B2(new_n356_), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT97), .B(KEYINPUT4), .Z(new_n386_));
  NAND4_X1  g185(.A1(new_n385_), .A2(new_n351_), .A3(new_n355_), .A4(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n348_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT98), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n348_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n396_));
  OR3_X1    g195(.A1(new_n388_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n394_), .B1(new_n388_), .B2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G227gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(G15gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n334_), .B(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n355_), .A2(new_n351_), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n405_), .B(KEYINPUT31), .Z(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(KEYINPUT81), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n308_), .B(new_n403_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n406_), .A2(KEYINPUT81), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G71gat), .B(G99gat), .ZN(new_n411_));
  INV_X1    g210(.A(G43gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(new_n410_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n400_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G228gat), .A2(G233gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT84), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n315_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n312_), .A2(new_n314_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n425_), .A2(new_n268_), .B1(new_n385_), .B2(KEYINPUT29), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n385_), .A2(KEYINPUT29), .ZN(new_n428_));
  INV_X1    g227(.A(new_n422_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n282_), .B(new_n428_), .C1(KEYINPUT84), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n421_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n282_), .A2(new_n428_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n282_), .A2(KEYINPUT84), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n422_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(new_n430_), .A3(new_n420_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT28), .B1(new_n385_), .B2(KEYINPUT29), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n365_), .A2(new_n376_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT28), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G22gat), .B(G50gat), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n438_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT88), .B1(new_n437_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n449_));
  AOI211_X1 g248(.A(new_n449_), .B(new_n446_), .C1(new_n432_), .C2(new_n436_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n420_), .B1(new_n435_), .B2(new_n430_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT90), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n446_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n436_), .A2(KEYINPUT89), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT89), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n435_), .A2(new_n455_), .A3(new_n430_), .A4(new_n420_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n452_), .B(new_n421_), .C1(new_n427_), .C2(new_n431_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  OAI22_X1  g257(.A1(new_n448_), .A2(new_n450_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n347_), .A2(new_n419_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n400_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n342_), .A2(new_n345_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n377_), .A2(new_n383_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n394_), .B1(new_n463_), .B2(new_n395_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n384_), .A2(new_n348_), .A3(new_n387_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT99), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n398_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n398_), .A2(new_n467_), .A3(KEYINPUT33), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n466_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(KEYINPUT32), .B(new_n205_), .C1(new_n318_), .C2(new_n323_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n336_), .A2(new_n340_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n474_), .A2(new_n475_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n462_), .A2(new_n472_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  OAI22_X1  g276(.A1(new_n461_), .A2(new_n347_), .B1(new_n477_), .B2(new_n459_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n417_), .A2(new_n418_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n460_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G29gat), .B(G36gat), .Z(new_n481_));
  XOR2_X1   g280(.A(G43gat), .B(G50gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486_));
  INV_X1    g285(.A(G1gat), .ZN(new_n487_));
  INV_X1    g286(.A(G8gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G8gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n490_), .B(new_n491_), .Z(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n485_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n483_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n492_), .A2(new_n483_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n495_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n496_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G113gat), .B(G141gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G169gat), .B(G197gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT74), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n502_), .B(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT101), .B1(new_n480_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT101), .ZN(new_n510_));
  INV_X1    g309(.A(new_n508_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n479_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n462_), .A2(new_n472_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n473_), .A2(new_n476_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n459_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n329_), .A2(new_n346_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n435_), .A2(new_n430_), .A3(new_n420_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n447_), .B1(new_n519_), .B2(new_n451_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n449_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n437_), .A2(KEYINPUT88), .A3(new_n447_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n453_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n452_), .A2(new_n451_), .B1(new_n436_), .B2(KEYINPUT89), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(new_n456_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n399_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n518_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n512_), .B1(new_n517_), .B2(new_n528_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n510_), .B(new_n511_), .C1(new_n529_), .C2(new_n460_), .ZN(new_n530_));
  INV_X1    g329(.A(G230gat), .ZN(new_n531_));
  INV_X1    g330(.A(G233gat), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G85gat), .ZN(new_n534_));
  INV_X1    g333(.A(G92gat), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT9), .ZN(new_n536_));
  XOR2_X1   g335(.A(G85gat), .B(G92gat), .Z(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(KEYINPUT9), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT10), .B(G99gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(G106gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT6), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n547_), .A2(KEYINPUT64), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(KEYINPUT64), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n544_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n538_), .A2(new_n542_), .A3(new_n546_), .A4(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT65), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT7), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n553_), .B(new_n554_), .C1(G99gat), .C2(G106gat), .ZN(new_n555_));
  INV_X1    g354(.A(G99gat), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n556_), .B(new_n541_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n550_), .A2(new_n546_), .A3(new_n552_), .A4(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT8), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n537_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n559_), .B2(new_n537_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n551_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G57gat), .B(G64gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT11), .ZN(new_n565_));
  XOR2_X1   g364(.A(G71gat), .B(G78gat), .Z(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n564_), .A2(KEYINPUT11), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n563_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n572_), .B(new_n551_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(KEYINPUT12), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n563_), .A2(new_n575_), .A3(new_n570_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n533_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT66), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n571_), .A2(new_n578_), .A3(new_n573_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n571_), .A2(new_n578_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n533_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n577_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G120gat), .B(G148gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  NOR2_X1   g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n582_), .A2(new_n579_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n574_), .A2(new_n576_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n581_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n592_), .A3(new_n588_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT68), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n583_), .A2(KEYINPUT68), .A3(new_n588_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n589_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n597_), .A2(KEYINPUT13), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(KEYINPUT13), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n509_), .A2(new_n530_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT73), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT16), .ZN(new_n604_));
  XOR2_X1   g403(.A(G183gat), .B(G211gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n602_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(new_n493_), .ZN(new_n609_));
  AND2_X1   g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n570_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n572_), .A3(new_n612_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n606_), .A2(new_n607_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n551_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n559_), .A2(new_n537_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT8), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n559_), .A2(new_n560_), .A3(new_n537_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT35), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT34), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n623_), .A2(new_n483_), .B1(new_n624_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n563_), .A2(new_n485_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(KEYINPUT70), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n627_), .A2(new_n624_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n628_), .B(new_n629_), .C1(KEYINPUT70), .C2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n633_), .A2(new_n635_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n633_), .A2(new_n635_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n638_), .B(KEYINPUT36), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT72), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT72), .ZN(new_n646_));
  AOI211_X1 g445(.A(new_n646_), .B(new_n643_), .C1(new_n633_), .C2(new_n635_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n641_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT37), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n642_), .A2(new_n644_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(KEYINPUT37), .A3(new_n641_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n601_), .A2(new_n618_), .A3(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n399_), .B(KEYINPUT102), .Z(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n487_), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n648_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT104), .B(new_n641_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n480_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n664_), .A2(new_n617_), .A3(new_n511_), .A4(new_n600_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G1gat), .B1(new_n665_), .B2(new_n400_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n658_), .A2(new_n659_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT105), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n658_), .A2(new_n669_), .A3(new_n659_), .A4(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1324gat));
  OAI21_X1  g470(.A(G8gat), .B1(new_n665_), .B2(new_n518_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT39), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n654_), .A2(new_n488_), .A3(new_n347_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n665_), .B2(new_n479_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT41), .Z(new_n679_));
  NAND3_X1  g478(.A1(new_n654_), .A2(new_n402_), .A3(new_n512_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1326gat));
  OAI21_X1  g480(.A(G22gat), .B1(new_n665_), .B2(new_n516_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT106), .Z(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT42), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(KEYINPUT42), .ZN(new_n685_));
  INV_X1    g484(.A(G22gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n654_), .A2(new_n686_), .A3(new_n459_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n685_), .A3(new_n687_), .ZN(G1327gat));
  INV_X1    g487(.A(new_n663_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n617_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n509_), .A2(new_n530_), .A3(new_n600_), .A4(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G29gat), .B1(new_n692_), .B2(new_n399_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n653_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n480_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n696_), .B(new_n653_), .C1(new_n529_), .C2(new_n460_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n600_), .A2(new_n618_), .A3(new_n511_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(KEYINPUT44), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n699_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n704_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n706_), .A2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n655_), .A2(G29gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n693_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n347_), .A2(new_n713_), .ZN(new_n714_));
  OR3_X1    g513(.A1(new_n691_), .A2(KEYINPUT45), .A3(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT45), .B1(new_n691_), .B2(new_n714_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n347_), .B1(new_n704_), .B2(KEYINPUT44), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n719_), .B2(new_n713_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n720_), .A2(KEYINPUT108), .A3(KEYINPUT46), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT46), .B1(new_n720_), .B2(KEYINPUT108), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  NOR2_X1   g522(.A1(new_n479_), .A2(new_n412_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n706_), .A2(new_n709_), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n412_), .B1(new_n691_), .B2(new_n479_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n692_), .B2(new_n459_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n459_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n710_), .B2(new_n730_), .ZN(G1331gat));
  NOR2_X1   g530(.A1(new_n600_), .A2(new_n511_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n664_), .A2(new_n732_), .A3(new_n617_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G57gat), .B1(new_n733_), .B2(new_n400_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n480_), .A2(new_n600_), .A3(new_n511_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n617_), .A3(new_n694_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n655_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(G57gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n736_), .B2(new_n738_), .ZN(G1332gat));
  OAI21_X1  g538(.A(G64gat), .B1(new_n733_), .B2(new_n518_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT48), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n518_), .A2(G64gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n736_), .B2(new_n742_), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n733_), .B2(new_n479_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT49), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n479_), .A2(G71gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n736_), .B2(new_n746_), .ZN(G1334gat));
  OAI21_X1  g546(.A(G78gat), .B1(new_n733_), .B2(new_n516_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT50), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n516_), .A2(G78gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n736_), .B2(new_n750_), .ZN(G1335gat));
  NAND2_X1  g550(.A1(new_n735_), .A2(new_n690_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT109), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n534_), .A3(new_n655_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n698_), .A2(new_n618_), .A3(new_n732_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT110), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(KEYINPUT110), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n400_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n758_), .B2(new_n534_), .ZN(G1336gat));
  NAND3_X1  g558(.A1(new_n753_), .A2(new_n535_), .A3(new_n347_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n756_), .A2(new_n757_), .A3(new_n518_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n535_), .ZN(G1337gat));
  OAI21_X1  g561(.A(G99gat), .B1(new_n755_), .B2(new_n479_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n753_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n512_), .A2(new_n540_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g566(.A(G106gat), .B1(new_n755_), .B2(new_n516_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT52), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT52), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n459_), .A2(new_n541_), .ZN(new_n771_));
  OAI22_X1  g570(.A1(new_n769_), .A2(new_n770_), .B1(new_n764_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  OAI221_X1 g573(.A(new_n774_), .B1(new_n764_), .B2(new_n771_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(G113gat), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n347_), .A2(new_n459_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n779_), .A2(new_n479_), .A3(new_n737_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n591_), .A2(KEYINPUT55), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n533_), .A2(KEYINPUT112), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n577_), .B2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n588_), .B1(new_n788_), .B2(new_n784_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n789_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n494_), .A2(new_n495_), .A3(new_n500_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n499_), .A2(new_n496_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n505_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n506_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT68), .B1(new_n583_), .B2(new_n588_), .ZN(new_n799_));
  AND4_X1   g598(.A1(KEYINPUT68), .A2(new_n590_), .A3(new_n592_), .A4(new_n588_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n782_), .B1(new_n792_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n787_), .A2(new_n789_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n789_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n797_), .B1(new_n596_), .B2(new_n595_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(KEYINPUT114), .A3(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n802_), .A2(new_n803_), .A3(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT115), .A3(new_n653_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(KEYINPUT58), .A3(new_n809_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT115), .B1(new_n811_), .B2(new_n653_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n799_), .A2(new_n800_), .B1(new_n583_), .B2(new_n588_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n508_), .B1(new_n596_), .B2(new_n595_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n820_), .A2(new_n798_), .B1(new_n808_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n819_), .B1(new_n822_), .B2(new_n663_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT57), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n819_), .B(new_n825_), .C1(new_n822_), .C2(new_n663_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n618_), .B1(new_n818_), .B2(new_n827_), .ZN(new_n828_));
  OR3_X1    g627(.A1(new_n618_), .A2(KEYINPUT111), .A3(new_n511_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT111), .B1(new_n618_), .B2(new_n511_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n600_), .A2(new_n694_), .A3(new_n829_), .A4(new_n830_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT54), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n781_), .B1(new_n828_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n777_), .B1(new_n834_), .B2(new_n508_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT59), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n811_), .A2(new_n653_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n824_), .A2(new_n826_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n617_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n831_), .B(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n780_), .B(new_n837_), .C1(new_n843_), .C2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n511_), .A2(G113gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT118), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n846_), .B(new_n848_), .C1(new_n833_), .C2(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n835_), .A2(new_n850_), .ZN(G1340gat));
  OAI21_X1  g650(.A(new_n846_), .B1(new_n833_), .B2(new_n849_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G120gat), .B1(new_n852_), .B2(new_n600_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G120gat), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n600_), .A2(KEYINPUT60), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n853_), .B1(new_n834_), .B2(new_n857_), .ZN(G1341gat));
  OAI21_X1  g657(.A(G127gat), .B1(new_n852_), .B2(new_n618_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n618_), .A2(G127gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n834_), .B2(new_n860_), .ZN(G1342gat));
  NAND2_X1  g660(.A1(new_n653_), .A2(G134gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT119), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n846_), .B(new_n863_), .C1(new_n833_), .C2(new_n849_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n663_), .B(new_n780_), .C1(new_n843_), .C2(new_n845_), .ZN(new_n865_));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n864_), .A2(KEYINPUT120), .A3(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1343gat));
  NOR2_X1   g671(.A1(new_n843_), .A2(new_n845_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n518_), .A2(new_n459_), .A3(new_n479_), .A4(new_n655_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT121), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n511_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g677(.A(new_n600_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n617_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  INV_X1    g683(.A(G162gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n876_), .A2(new_n885_), .A3(new_n663_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n876_), .A2(new_n653_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n886_), .B1(new_n888_), .B2(new_n885_), .ZN(G1347gat));
  NOR4_X1   g688(.A1(new_n518_), .A2(new_n655_), .A3(new_n459_), .A4(new_n479_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n511_), .B(new_n890_), .C1(new_n843_), .C2(new_n845_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT122), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n828_), .A2(new_n832_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n893_), .A2(new_n894_), .A3(new_n511_), .A4(new_n890_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(new_n895_), .A3(G169gat), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n892_), .A2(new_n895_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n893_), .A2(new_n890_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(new_n216_), .A3(new_n511_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n899_), .A3(new_n901_), .ZN(G1348gat));
  NAND3_X1  g701(.A1(new_n893_), .A2(new_n879_), .A3(new_n890_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(KEYINPUT123), .B2(new_n217_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n217_), .A2(KEYINPUT123), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT124), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n904_), .B(new_n906_), .ZN(G1349gat));
  NAND2_X1  g706(.A1(new_n900_), .A2(new_n617_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n234_), .ZN(new_n909_));
  AOI21_X1  g708(.A(G183gat), .B1(new_n900_), .B2(new_n617_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1350gat));
  NAND2_X1  g710(.A1(new_n900_), .A2(new_n653_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G190gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n663_), .A2(new_n235_), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT125), .Z(new_n915_));
  NAND2_X1  g714(.A1(new_n900_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n916_), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n527_), .A2(new_n347_), .A3(new_n479_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n873_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n511_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n879_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n275_), .A2(KEYINPUT126), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n275_), .A2(KEYINPUT126), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n922_), .B2(new_n923_), .ZN(G1353gat));
  XOR2_X1   g725(.A(KEYINPUT63), .B(G211gat), .Z(new_n927_));
  AND3_X1   g726(.A1(new_n919_), .A2(new_n617_), .A3(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n919_), .A2(new_n617_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n928_), .B1(new_n929_), .B2(new_n930_), .ZN(G1354gat));
  AOI21_X1  g730(.A(G218gat), .B1(new_n919_), .B2(new_n663_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n653_), .A2(G218gat), .ZN(new_n933_));
  XOR2_X1   g732(.A(new_n933_), .B(KEYINPUT127), .Z(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n919_), .B2(new_n934_), .ZN(G1355gat));
endmodule


