//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT81), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT81), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(G169gat), .B2(G176gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n203_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT83), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n214_), .B(KEYINPUT82), .Z(new_n215_));
  NAND2_X1  g014(.A1(new_n206_), .A2(new_n208_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n203_), .A2(new_n210_), .A3(KEYINPUT83), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT79), .B(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT26), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT80), .B1(new_n222_), .B2(KEYINPUT26), .ZN(new_n223_));
  OR3_X1    g022(.A1(new_n222_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n220_), .A2(new_n221_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n213_), .A2(new_n217_), .A3(new_n218_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G169gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n204_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n205_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT85), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(new_n202_), .B2(KEYINPUT23), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n232_), .B1(new_n203_), .B2(new_n231_), .ZN(new_n233_));
  INV_X1    g032(.A(G183gat), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n219_), .A2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n230_), .B(new_n215_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n226_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT30), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G43gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n237_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G43gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G15gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G71gat), .B(G99gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  NAND3_X1  g046(.A1(new_n239_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n239_), .B2(new_n243_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT86), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G113gat), .ZN(new_n254_));
  INV_X1    g053(.A(G127gat), .ZN(new_n255_));
  INV_X1    g054(.A(G134gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G113gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G127gat), .A2(G134gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n254_), .A2(new_n260_), .A3(G120gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(G120gat), .B1(new_n254_), .B2(new_n260_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT31), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n252_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n250_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT86), .B1(new_n266_), .B2(new_n248_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n264_), .B1(new_n267_), .B2(new_n252_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G1gat), .B(G29gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G57gat), .B(G85gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT88), .B(KEYINPUT3), .ZN(new_n276_));
  OR2_X1    g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT89), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT89), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n281_), .A2(KEYINPUT88), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(KEYINPUT88), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n279_), .B(new_n280_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT2), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT2), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(G141gat), .A3(G148gat), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n286_), .A2(new_n288_), .B1(new_n277_), .B2(KEYINPUT3), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n278_), .A2(new_n284_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G155gat), .ZN(new_n291_));
  INV_X1    g090(.A(G162gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(KEYINPUT87), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT87), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(G155gat), .B2(G162gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n290_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n296_), .B(KEYINPUT1), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n293_), .A2(new_n295_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n277_), .B(new_n285_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n261_), .A2(new_n262_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(new_n303_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n263_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(KEYINPUT96), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT96), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n263_), .A2(new_n298_), .A3(new_n312_), .A4(new_n301_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n308_), .B1(new_n314_), .B2(KEYINPUT4), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n307_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n275_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n306_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n304_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n318_), .B(new_n274_), .C1(new_n319_), .C2(new_n308_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(KEYINPUT101), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(KEYINPUT4), .ZN(new_n322_));
  INV_X1    g121(.A(new_n308_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT101), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(new_n318_), .A4(new_n274_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n269_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT93), .ZN(new_n331_));
  INV_X1    g130(.A(G197gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT91), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT91), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(G197gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n331_), .B1(new_n336_), .B2(G204gat), .ZN(new_n337_));
  INV_X1    g136(.A(G204gat), .ZN(new_n338_));
  AOI211_X1 g137(.A(KEYINPUT93), .B(new_n338_), .C1(new_n333_), .C2(new_n335_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT94), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT21), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT92), .B1(new_n332_), .B2(G204gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT92), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(new_n338_), .A3(G197gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .A4(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G211gat), .B(G218gat), .Z(new_n348_));
  NOR2_X1   g147(.A1(new_n332_), .A2(new_n338_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n350_), .B2(KEYINPUT21), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT91), .B(G197gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT93), .B1(new_n352_), .B2(new_n338_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n334_), .A2(G197gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n332_), .A2(KEYINPUT91), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n331_), .B(G204gat), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n353_), .A2(new_n342_), .A3(new_n356_), .A4(new_n346_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT94), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n347_), .A2(new_n351_), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n353_), .A2(new_n356_), .A3(new_n346_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(KEYINPUT21), .A3(new_n348_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT26), .B(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n221_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT95), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n233_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n363_), .A2(KEYINPUT95), .A3(new_n365_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT22), .B(G169gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n205_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n215_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n362_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT19), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n226_), .A2(new_n236_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n378_), .A2(KEYINPUT20), .A3(new_n381_), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT100), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT20), .ZN(new_n386_));
  INV_X1    g185(.A(new_n361_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n357_), .B(new_n341_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n351_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n389_), .B2(new_n382_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT100), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n381_), .A4(new_n378_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n362_), .A2(new_n237_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT20), .B1(new_n362_), .B2(new_n377_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n380_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n385_), .A2(new_n392_), .A3(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT18), .B(G64gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(G92gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n397_), .A2(KEYINPUT103), .A3(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n403_), .A2(KEYINPUT27), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(new_n402_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT103), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n381_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n390_), .A2(new_n378_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n407_), .B1(new_n381_), .B2(new_n408_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n405_), .A2(new_n406_), .B1(new_n409_), .B2(new_n401_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT27), .ZN(new_n411_));
  INV_X1    g210(.A(new_n377_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n386_), .B1(new_n389_), .B2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n380_), .B1(new_n413_), .B2(new_n393_), .ZN(new_n414_));
  AND4_X1   g213(.A1(KEYINPUT20), .A2(new_n378_), .A3(new_n380_), .A4(new_n383_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n401_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n407_), .B(new_n402_), .C1(new_n381_), .C2(new_n408_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n404_), .A2(new_n410_), .B1(new_n411_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT104), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n302_), .A2(KEYINPUT29), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n362_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n423_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G228gat), .A2(G233gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n424_), .A2(G228gat), .A3(G233gat), .A4(new_n425_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(KEYINPUT90), .A3(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n302_), .A2(KEYINPUT29), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT28), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G22gat), .B(G50gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n430_), .B(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n419_), .A2(new_n420_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n420_), .B1(new_n419_), .B2(new_n435_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n330_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n401_), .A2(KEYINPUT32), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n409_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n439_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n397_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n327_), .A2(KEYINPUT102), .A3(new_n440_), .A4(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n442_), .A2(new_n440_), .A3(new_n321_), .A4(new_n326_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT102), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n320_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT98), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n320_), .A2(KEYINPUT98), .A3(new_n448_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n324_), .A2(KEYINPUT33), .A3(new_n318_), .A4(new_n274_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n416_), .A2(new_n417_), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n322_), .A2(new_n306_), .A3(new_n305_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n314_), .A2(new_n307_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n275_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(new_n455_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT99), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT99), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n453_), .A2(new_n455_), .A3(new_n461_), .A4(new_n458_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n447_), .A2(new_n435_), .A3(new_n460_), .A4(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n405_), .A2(new_n406_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n464_), .A2(KEYINPUT27), .A3(new_n416_), .A4(new_n403_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n418_), .A2(new_n411_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n328_), .A3(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n430_), .B(new_n434_), .Z(new_n468_));
  AOI21_X1  g267(.A(new_n269_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n463_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n438_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G50gat), .ZN(new_n472_));
  INV_X1    g271(.A(G29gat), .ZN(new_n473_));
  INV_X1    g272(.A(G36gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G29gat), .A2(G36gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n242_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n242_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n472_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n479_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G50gat), .A3(new_n477_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n480_), .A2(new_n482_), .A3(KEYINPUT15), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT15), .B1(new_n480_), .B2(new_n482_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G15gat), .B(G22gat), .Z(new_n487_));
  NAND2_X1  g286(.A1(G1gat), .A2(G8gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n487_), .B1(KEYINPUT14), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT76), .ZN(new_n490_));
  XOR2_X1   g289(.A(G1gat), .B(G8gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  MUX2_X1   g291(.A(new_n483_), .B(new_n486_), .S(new_n492_), .Z(new_n493_));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n492_), .B(new_n483_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n494_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT78), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G113gat), .B(G141gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(G197gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT77), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(new_n204_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n501_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G57gat), .B(G64gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT67), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT11), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G71gat), .B(G78gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT11), .ZN(new_n514_));
  OR3_X1    g313(.A1(new_n509_), .A2(new_n514_), .A3(new_n512_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G85gat), .B(G92gat), .Z(new_n516_));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n519_), .B(new_n520_), .C1(new_n521_), .C2(KEYINPUT7), .ZN(new_n522_));
  INV_X1    g321(.A(G99gat), .ZN(new_n523_));
  INV_X1    g322(.A(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n523_), .B(new_n524_), .C1(new_n525_), .C2(KEYINPUT66), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n521_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n516_), .B1(new_n522_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT8), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT8), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n531_), .B(new_n516_), .C1(new_n522_), .C2(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n519_), .A2(new_n520_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n516_), .B2(KEYINPUT9), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT64), .ZN(new_n536_));
  INV_X1    g335(.A(G92gat), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT9), .ZN(new_n538_));
  NOR2_X1   g337(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(G85gat), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT10), .B(G99gat), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n524_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n535_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT65), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n535_), .A2(KEYINPUT65), .A3(new_n540_), .A4(new_n542_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n533_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n513_), .A2(new_n515_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n513_), .A2(new_n515_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n547_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n555_), .A2(new_n556_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n552_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n548_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n553_), .A2(new_n554_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(new_n556_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n548_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(G230gat), .A3(G233gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(G120gat), .B(G148gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  NAND3_X1  g367(.A1(new_n560_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT70), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n560_), .A2(new_n563_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n568_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT13), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(KEYINPUT13), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n507_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n471_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n555_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n492_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT16), .B(G183gat), .ZN(new_n583_));
  INV_X1    g382(.A(G211gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n582_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n587_), .A2(new_n588_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(new_n582_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(G134gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n292_), .ZN(new_n597_));
  INV_X1    g396(.A(G232gat), .ZN(new_n598_));
  INV_X1    g397(.A(G233gat), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n486_), .A2(new_n547_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n533_), .A2(new_n545_), .A3(new_n546_), .A4(new_n483_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT72), .Z(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n601_), .A2(new_n602_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n600_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(KEYINPUT73), .A3(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n605_), .A2(new_n608_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n609_), .B2(KEYINPUT73), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n604_), .B(new_n600_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n607_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT35), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n612_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n603_), .A2(KEYINPUT35), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n594_), .B(new_n597_), .C1(new_n617_), .C2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n608_), .B1(new_n605_), .B2(new_n611_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n613_), .A2(new_n614_), .A3(new_n607_), .ZN(new_n622_));
  OAI22_X1  g421(.A1(new_n621_), .A2(new_n622_), .B1(KEYINPUT35), .B2(new_n603_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n597_), .A2(new_n594_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n597_), .A2(new_n594_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n612_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .A4(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n620_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT37), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT74), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(KEYINPUT74), .A3(KEYINPUT37), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT75), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n628_), .B2(KEYINPUT37), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT37), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n620_), .A2(new_n627_), .A3(KEYINPUT75), .A4(new_n635_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n631_), .A2(new_n632_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n578_), .A2(new_n593_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(G1gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n327_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT38), .ZN(new_n641_));
  INV_X1    g440(.A(new_n628_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n578_), .A2(new_n593_), .A3(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(new_n327_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n641_), .B1(new_n639_), .B2(new_n644_), .ZN(G1324gat));
  NAND2_X1  g444(.A1(new_n465_), .A2(new_n466_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G8gat), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(KEYINPUT39), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(G8gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n638_), .A2(new_n653_), .A3(new_n646_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n648_), .A2(new_n649_), .A3(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n652_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g457(.A(G15gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n643_), .B2(new_n269_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT41), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n638_), .A2(new_n659_), .A3(new_n269_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1326gat));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n643_), .B2(new_n468_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT42), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n638_), .A2(new_n664_), .A3(new_n468_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1327gat));
  OR3_X1    g467(.A1(new_n628_), .A2(KEYINPUT108), .A3(new_n592_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT108), .B1(new_n628_), .B2(new_n592_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n463_), .A2(new_n469_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n646_), .B2(new_n468_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n419_), .A2(new_n420_), .A3(new_n435_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n329_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n577_), .B(new_n671_), .C1(new_n672_), .C2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT109), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n471_), .A2(new_n678_), .A3(new_n577_), .A4(new_n671_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n327_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n637_), .C1(new_n672_), .C2(new_n675_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n673_), .A2(new_n674_), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n686_), .A2(new_n330_), .B1(new_n463_), .B2(new_n469_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n637_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n471_), .A2(KEYINPUT106), .A3(new_n682_), .A4(new_n637_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n685_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n577_), .A2(new_n593_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(KEYINPUT44), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n691_), .A2(new_n693_), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n473_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n681_), .B1(new_n699_), .B2(new_n327_), .ZN(G1328gat));
  NOR2_X1   g499(.A1(new_n697_), .A2(new_n698_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n474_), .B1(new_n701_), .B2(new_n646_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n677_), .A2(new_n474_), .A3(new_n646_), .A4(new_n679_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(KEYINPUT110), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(KEYINPUT110), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n680_), .A2(new_n708_), .A3(new_n474_), .A4(new_n646_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n704_), .A2(KEYINPUT110), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(KEYINPUT45), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT111), .B1(new_n702_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n691_), .A2(new_n693_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n695_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n691_), .A2(new_n693_), .A3(new_n696_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n646_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n711_), .A4(new_n707_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n713_), .A2(KEYINPUT46), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT46), .B1(new_n713_), .B2(new_n720_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  AND3_X1   g522(.A1(new_n680_), .A2(new_n242_), .A3(new_n269_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n701_), .A2(new_n269_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(G43gat), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n680_), .B2(new_n468_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n697_), .A2(new_n698_), .A3(new_n435_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G50gat), .ZN(G1331gat));
  NAND2_X1  g529(.A1(new_n575_), .A2(new_n576_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(new_n506_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n471_), .A2(new_n732_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n733_), .A2(new_n592_), .A3(new_n628_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(G57gat), .A3(new_n327_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n637_), .A2(new_n593_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n737_), .A2(new_n328_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(G57gat), .B2(new_n738_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT112), .Z(G1332gat));
  INV_X1    g539(.A(G64gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n734_), .B2(new_n646_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT48), .Z(new_n743_));
  INV_X1    g542(.A(new_n737_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(new_n741_), .A3(new_n646_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n734_), .B2(new_n269_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT113), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT49), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n744_), .A2(new_n747_), .A3(new_n269_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n734_), .B2(new_n468_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT50), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n744_), .A2(new_n753_), .A3(new_n468_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n733_), .A2(new_n671_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT114), .ZN(new_n759_));
  AOI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n327_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n732_), .A2(new_n593_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT115), .Z(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(new_n691_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n763_), .A2(G85gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n760_), .B1(new_n327_), .B2(new_n764_), .ZN(G1336gat));
  AOI21_X1  g564(.A(G92gat), .B1(new_n759_), .B2(new_n646_), .ZN(new_n766_));
  XOR2_X1   g565(.A(KEYINPUT64), .B(G92gat), .Z(new_n767_));
  NOR2_X1   g566(.A1(new_n419_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n763_), .B2(new_n768_), .ZN(G1337gat));
  NAND3_X1  g568(.A1(new_n759_), .A2(new_n541_), .A3(new_n269_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n763_), .A2(new_n269_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n523_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n762_), .A2(new_n691_), .A3(new_n468_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G106gat), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT116), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n777_), .A3(G106gat), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n759_), .A2(new_n524_), .A3(new_n468_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n776_), .A2(KEYINPUT52), .A3(new_n778_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n781_), .A2(new_n785_), .A3(new_n782_), .A4(new_n783_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1339gat));
  NAND3_X1  g588(.A1(new_n686_), .A2(new_n327_), .A3(new_n269_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT122), .ZN(new_n791_));
  NOR2_X1   g590(.A1(KEYINPUT118), .A2(KEYINPUT55), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n560_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n553_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(G230gat), .A3(G233gat), .ZN(new_n795_));
  AND2_X1   g594(.A1(KEYINPUT118), .A2(KEYINPUT55), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n560_), .B1(new_n792_), .B2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n793_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT119), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n793_), .A2(new_n795_), .A3(new_n797_), .A4(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n799_), .A2(new_n800_), .A3(new_n572_), .A4(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(new_n570_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n495_), .A2(new_n498_), .A3(new_n505_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n493_), .A2(new_n494_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n496_), .A2(new_n497_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n805_), .B1(new_n505_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n799_), .A2(new_n572_), .A3(new_n802_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(KEYINPUT56), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT121), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n804_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n814_), .B1(new_n804_), .B2(new_n811_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n791_), .B1(new_n818_), .B2(new_n688_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n809_), .B1(new_n573_), .B2(new_n570_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n810_), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n821_), .A2(new_n506_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n570_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n810_), .A2(KEYINPUT120), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n800_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n820_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  OR3_X1    g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n642_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n826_), .B2(new_n642_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n817_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n815_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(KEYINPUT122), .A3(new_n637_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n819_), .A2(new_n828_), .A3(new_n829_), .A4(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n593_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n688_), .A2(new_n592_), .A3(new_n507_), .A4(new_n731_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT54), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n790_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837_), .B2(new_n506_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n831_), .A2(new_n637_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n828_), .A2(new_n829_), .A3(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n836_), .B1(new_n840_), .B2(new_n592_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n837_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n258_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n838_), .B1(new_n846_), .B2(new_n506_), .ZN(G1340gat));
  OAI21_X1  g646(.A(G120gat), .B1(new_n845_), .B2(new_n731_), .ZN(new_n848_));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n731_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n837_), .B(new_n850_), .C1(KEYINPUT60), .C2(new_n849_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(G1341gat));
  OAI211_X1 g651(.A(new_n843_), .B(new_n592_), .C1(new_n837_), .C2(new_n844_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G127gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n837_), .A2(new_n255_), .A3(new_n592_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT123), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n854_), .A2(new_n858_), .A3(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1342gat));
  AOI21_X1  g659(.A(G134gat), .B1(new_n837_), .B2(new_n642_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n845_), .A2(new_n256_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n637_), .ZN(G1343gat));
  NAND2_X1  g662(.A1(new_n834_), .A2(new_n836_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n269_), .A2(new_n435_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n419_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n865_), .A2(new_n328_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n506_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g669(.A(new_n731_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g672(.A1(new_n868_), .A2(new_n592_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  AOI21_X1  g675(.A(G162gat), .B1(new_n868_), .B2(new_n642_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n637_), .A2(G162gat), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT124), .Z(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n868_), .B2(new_n879_), .ZN(G1347gat));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n329_), .A2(new_n419_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n841_), .A2(new_n435_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n506_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n881_), .B1(new_n885_), .B2(G169gat), .ZN(new_n886_));
  AOI211_X1 g685(.A(KEYINPUT62), .B(new_n204_), .C1(new_n884_), .C2(new_n506_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n506_), .A2(new_n374_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(KEYINPUT125), .Z(new_n889_));
  OAI22_X1  g688(.A1(new_n886_), .A2(new_n887_), .B1(new_n883_), .B2(new_n889_), .ZN(G1348gat));
  AOI21_X1  g689(.A(G176gat), .B1(new_n884_), .B2(new_n871_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n864_), .A2(new_n435_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n892_), .A2(new_n205_), .A3(new_n731_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n882_), .B2(new_n893_), .ZN(G1349gat));
  NOR3_X1   g693(.A1(new_n883_), .A2(new_n593_), .A3(new_n221_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n895_), .A2(KEYINPUT126), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n882_), .A2(new_n592_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n234_), .B1(new_n892_), .B2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n895_), .A2(KEYINPUT126), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n896_), .A2(new_n898_), .A3(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n883_), .B2(new_n688_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n642_), .A2(new_n364_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n883_), .B2(new_n902_), .ZN(G1351gat));
  AND2_X1   g702(.A1(new_n864_), .A2(new_n866_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n419_), .A2(new_n327_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(new_n506_), .A3(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g706(.A1(new_n904_), .A2(new_n871_), .A3(new_n905_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G204gat), .ZN(G1353gat));
  AND4_X1   g708(.A1(new_n592_), .A2(new_n864_), .A3(new_n866_), .A4(new_n905_), .ZN(new_n910_));
  OR2_X1    g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  OR3_X1    g710(.A1(new_n910_), .A2(KEYINPUT127), .A3(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT127), .B1(new_n910_), .B2(new_n911_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT63), .B(G211gat), .Z(new_n914_));
  AOI22_X1  g713(.A1(new_n912_), .A2(new_n913_), .B1(new_n910_), .B2(new_n914_), .ZN(G1354gat));
  AND3_X1   g714(.A1(new_n904_), .A2(G218gat), .A3(new_n905_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n904_), .A2(new_n642_), .A3(new_n905_), .ZN(new_n917_));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n916_), .A2(new_n637_), .B1(new_n917_), .B2(new_n918_), .ZN(G1355gat));
endmodule


