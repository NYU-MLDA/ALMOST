//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  OAI22_X1  g004(.A1(new_n203_), .A2(new_n204_), .B1(new_n205_), .B2(KEYINPUT94), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n204_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT95), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(KEYINPUT95), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n206_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n205_), .A2(KEYINPUT94), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n211_), .B(new_n212_), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n217_), .B(KEYINPUT96), .Z(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(KEYINPUT1), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n215_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT92), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n215_), .A3(KEYINPUT92), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n223_), .B(new_n224_), .C1(KEYINPUT1), .C2(new_n216_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT93), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n211_), .A2(new_n203_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n225_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n226_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n219_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G113gat), .B(G120gat), .ZN(new_n232_));
  INV_X1    g031(.A(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT91), .B(G127gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n202_), .B1(new_n231_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n202_), .A3(new_n237_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n225_), .A2(new_n228_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT93), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n225_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n243_), .A2(new_n244_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT103), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n236_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT103), .B1(new_n231_), .B2(new_n237_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n241_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT4), .B1(new_n231_), .B2(new_n237_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n240_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n248_), .B(new_n247_), .C1(new_n253_), .C2(new_n238_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n254_), .B2(KEYINPUT4), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n255_), .B2(new_n250_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G1gat), .B(G29gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G85gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT0), .B(G57gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n251_), .B(new_n260_), .C1(new_n255_), .C2(new_n250_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G197gat), .B(G204gat), .Z(new_n266_));
  AND3_X1   g065(.A1(new_n266_), .A2(KEYINPUT98), .A3(KEYINPUT21), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(KEYINPUT21), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G211gat), .B(G218gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  OR3_X1    g069(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n270_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(new_n231_), .B2(KEYINPUT29), .ZN(new_n274_));
  AND2_X1   g073(.A1(G228gat), .A2(G233gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n276_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G78gat), .B(G106gat), .Z(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n274_), .A2(new_n276_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n282_), .B1(new_n283_), .B2(new_n277_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n283_), .A2(new_n277_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT99), .B1(new_n286_), .B2(new_n280_), .ZN(new_n287_));
  XOR2_X1   g086(.A(KEYINPUT97), .B(KEYINPUT28), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n245_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G22gat), .B(G50gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n231_), .A2(KEYINPUT29), .ZN(new_n294_));
  INV_X1    g093(.A(new_n292_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n289_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n292_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n295_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(new_n288_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n285_), .B1(new_n287_), .B2(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n297_), .A2(new_n300_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n303_), .A2(KEYINPUT99), .A3(new_n281_), .A4(new_n284_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT20), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT25), .B(G183gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G190gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT82), .ZN(new_n310_));
  INV_X1    g109(.A(G190gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT26), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT82), .B1(new_n308_), .B2(G190gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n307_), .A2(new_n309_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT83), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G169gat), .ZN(new_n317_));
  INV_X1    g116(.A(G176gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(KEYINPUT24), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n321_));
  INV_X1    g120(.A(G183gat), .ZN(new_n322_));
  OR3_X1    g121(.A1(new_n322_), .A2(new_n311_), .A3(KEYINPUT23), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT23), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(KEYINPUT24), .A3(new_n319_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n316_), .A2(new_n321_), .A3(new_n326_), .A4(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT85), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT22), .B1(new_n332_), .B2(new_n317_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT22), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(KEYINPUT85), .A3(G169gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n318_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n329_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT86), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n324_), .A2(KEYINPUT87), .A3(KEYINPUT23), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT87), .B1(new_n324_), .B2(KEYINPUT23), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n323_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n336_), .A2(new_n329_), .A3(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n338_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n331_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT88), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n331_), .A2(new_n347_), .A3(KEYINPUT88), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n271_), .A2(new_n272_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n306_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT101), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT19), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n311_), .A2(KEYINPUT26), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n307_), .A2(new_n359_), .A3(new_n309_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n319_), .A2(KEYINPUT24), .A3(new_n327_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n320_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n341_), .A2(new_n360_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT100), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n326_), .A2(new_n343_), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT22), .B(G169gat), .Z(new_n367_));
  OAI211_X1 g166(.A(new_n366_), .B(new_n329_), .C1(G176gat), .C2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n273_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n354_), .A2(new_n355_), .A3(new_n358_), .A4(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n365_), .A2(new_n368_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n353_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n372_), .B(KEYINPUT20), .C1(new_n352_), .C2(new_n353_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n357_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n331_), .A2(KEYINPUT88), .A3(new_n347_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT88), .B1(new_n331_), .B2(new_n347_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n353_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n377_), .A2(KEYINPUT20), .A3(new_n369_), .A4(new_n358_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT101), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n370_), .A2(new_n374_), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381_));
  INV_X1    g180(.A(G92gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT18), .B(G64gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387_));
  INV_X1    g186(.A(new_n385_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n370_), .A2(new_n374_), .A3(new_n379_), .A4(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n273_), .A2(new_n368_), .A3(new_n363_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n354_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT106), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n357_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n377_), .A2(KEYINPUT20), .A3(new_n391_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT106), .B1(new_n395_), .B2(new_n358_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n373_), .A2(new_n357_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n394_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n385_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n370_), .A2(new_n379_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n400_), .A2(KEYINPUT107), .A3(new_n388_), .A4(new_n374_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT107), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n389_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n390_), .B1(new_n404_), .B2(KEYINPUT27), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n305_), .B1(new_n405_), .B2(new_n264_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n263_), .A2(KEYINPUT33), .ZN(new_n407_));
  INV_X1    g206(.A(new_n250_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(new_n241_), .B2(new_n249_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n410_), .B2(new_n252_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n251_), .A4(new_n260_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n386_), .A2(new_n389_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n250_), .B1(new_n410_), .B2(new_n252_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n241_), .A2(new_n249_), .A3(new_n408_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n261_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT104), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n416_), .A2(KEYINPUT104), .A3(new_n261_), .A4(new_n417_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n414_), .A2(new_n415_), .A3(new_n420_), .A4(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT105), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n388_), .A2(KEYINPUT32), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n380_), .B2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n380_), .A2(new_n424_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n424_), .B2(new_n398_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n264_), .B(new_n425_), .C1(new_n427_), .C2(new_n423_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n305_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n422_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT30), .B1(new_n375_), .B2(new_n376_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT30), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n350_), .A2(new_n432_), .A3(new_n351_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT90), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT31), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G227gat), .A2(G233gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT89), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G15gat), .B(G43gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G71gat), .B(G99gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n435_), .A2(new_n436_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT90), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n442_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT31), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n237_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n434_), .A2(KEYINPUT90), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n443_), .A2(new_n447_), .A3(new_n237_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n443_), .A2(new_n447_), .A3(new_n237_), .ZN(new_n453_));
  OAI22_X1  g252(.A1(new_n453_), .A2(new_n448_), .B1(KEYINPUT90), .B2(new_n434_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n406_), .A2(new_n430_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n305_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n389_), .B(KEYINPUT107), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n387_), .B1(new_n458_), .B2(new_n399_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n457_), .B(new_n265_), .C1(new_n459_), .C2(new_n390_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT108), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n404_), .A2(KEYINPUT27), .ZN(new_n463_));
  INV_X1    g262(.A(new_n390_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n264_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT108), .B1(new_n465_), .B2(new_n457_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n456_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G230gat), .A2(G233gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n468_), .B(KEYINPUT64), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT12), .ZN(new_n471_));
  INV_X1    g270(.A(G99gat), .ZN(new_n472_));
  INV_X1    g271(.A(G106gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT6), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(G99gat), .A3(G106gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT9), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(G85gat), .A3(G92gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G85gat), .B(G92gat), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n477_), .B(new_n479_), .C1(new_n478_), .C2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT10), .B(G99gat), .Z(new_n482_));
  AND2_X1   g281(.A1(new_n482_), .A2(new_n473_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT7), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n485_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n472_), .A2(new_n473_), .ZN(new_n491_));
  AND2_X1   g290(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT69), .B1(new_n490_), .B2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n474_), .A2(new_n476_), .A3(KEYINPUT68), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT68), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n477_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n491_), .B1(new_n492_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT69), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n485_), .A2(new_n489_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .A4(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n480_), .B(KEYINPUT67), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT70), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n503_), .A2(KEYINPUT70), .A3(new_n504_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(KEYINPUT8), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n477_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n510_), .A2(KEYINPUT66), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT8), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(KEYINPUT66), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n504_), .A4(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n484_), .B1(new_n509_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G57gat), .B(G64gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT11), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G71gat), .B(G78gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n516_), .B(KEYINPUT11), .Z(new_n520_));
  OAI21_X1  g319(.A(new_n519_), .B1(new_n520_), .B2(new_n518_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n471_), .B1(new_n515_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n484_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n503_), .A2(KEYINPUT70), .A3(new_n504_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT70), .B1(new_n503_), .B2(new_n504_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n512_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n514_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n521_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n523_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n471_), .A3(new_n521_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n470_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT5), .B(G176gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G204gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(G120gat), .B(G148gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT72), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n515_), .A2(new_n522_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT71), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n529_), .B2(new_n521_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n541_), .B(new_n470_), .C1(new_n543_), .C2(new_n540_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n534_), .A2(new_n539_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n539_), .B1(new_n534_), .B2(new_n544_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT13), .ZN(new_n547_));
  OR3_X1    g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G15gat), .B(G22gat), .Z(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT75), .B(G8gat), .Z(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(G1gat), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n551_), .B1(new_n553_), .B2(KEYINPUT14), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT76), .B(KEYINPUT77), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G1gat), .B(G8gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n556_), .B(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G43gat), .B(G50gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(G29gat), .B(G36gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT79), .B1(new_n559_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n559_), .B2(new_n563_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n556_), .B(new_n557_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(KEYINPUT79), .A3(new_n562_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n565_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n562_), .B(KEYINPUT15), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n559_), .A2(KEYINPUT80), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n559_), .A2(new_n563_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT80), .B1(new_n559_), .B2(new_n571_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n572_), .A2(new_n566_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT81), .B(G113gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G141gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G169gat), .B(G197gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n570_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n550_), .A2(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n467_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n515_), .B2(new_n571_), .ZN(new_n596_));
  AOI211_X1 g395(.A(new_n484_), .B(new_n562_), .C1(new_n509_), .C2(new_n514_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT73), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n571_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n529_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n515_), .A2(new_n563_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT73), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .A4(new_n595_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n593_), .A2(new_n594_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n598_), .A2(new_n605_), .A3(new_n603_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n590_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n590_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n608_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT74), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n609_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT74), .B1(new_n607_), .B2(new_n608_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT36), .B1(new_n616_), .B2(new_n610_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT37), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n598_), .A2(new_n605_), .A3(new_n603_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n605_), .B1(new_n598_), .B2(new_n603_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n612_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n614_), .A3(new_n590_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n609_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n617_), .A2(KEYINPUT37), .A3(new_n622_), .A4(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n618_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n559_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(new_n522_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G127gat), .B(G155gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(G211gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(KEYINPUT16), .B(G183gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(KEYINPUT17), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n629_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT78), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n633_), .A2(KEYINPUT17), .ZN(new_n637_));
  OR3_X1    g436(.A1(new_n629_), .A2(new_n634_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n626_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n587_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT109), .ZN(new_n642_));
  INV_X1    g441(.A(new_n640_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n467_), .A2(new_n586_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT109), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI211_X1 g446(.A(G1gat), .B(new_n265_), .C1(new_n642_), .C2(new_n647_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(KEYINPUT38), .ZN(new_n649_));
  INV_X1    g448(.A(new_n617_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n622_), .A2(new_n623_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n639_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n587_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G1gat), .B1(new_n655_), .B2(new_n265_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n648_), .A2(KEYINPUT38), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n649_), .A2(new_n656_), .A3(new_n657_), .ZN(G1324gat));
  NAND3_X1  g457(.A1(new_n587_), .A2(new_n654_), .A3(new_n405_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  AND4_X1   g459(.A1(KEYINPUT110), .A2(new_n659_), .A3(new_n660_), .A4(G8gat), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(KEYINPUT110), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n659_), .A2(G8gat), .B1(KEYINPUT110), .B2(new_n660_), .ZN(new_n663_));
  OR3_X1    g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n552_), .B1(new_n642_), .B2(new_n647_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n405_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n664_), .A2(KEYINPUT40), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n665_), .A2(new_n405_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n668_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n667_), .A2(new_n671_), .ZN(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n655_), .B2(new_n455_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT41), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n641_), .A2(G15gat), .A3(new_n455_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1326gat));
  OAI21_X1  g475(.A(G22gat), .B1(new_n655_), .B2(new_n429_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n429_), .A2(G22gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n641_), .B2(new_n679_), .ZN(G1327gat));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT37), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n624_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n683_), .A2(KEYINPUT111), .A3(new_n624_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n467_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n460_), .A2(new_n461_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n465_), .A2(KEYINPUT108), .A3(new_n457_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT43), .B1(new_n691_), .B2(new_n456_), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n688_), .A2(KEYINPUT43), .B1(new_n692_), .B2(new_n626_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n586_), .A2(new_n639_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n681_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n694_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  INV_X1    g496(.A(new_n687_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT111), .B1(new_n683_), .B2(new_n624_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n700_), .B2(new_n467_), .ZN(new_n701_));
  AOI211_X1 g500(.A(KEYINPUT43), .B(new_n684_), .C1(new_n691_), .C2(new_n456_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT44), .B(new_n696_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n695_), .A2(new_n703_), .A3(new_n264_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G29gat), .ZN(new_n705_));
  INV_X1    g504(.A(new_n639_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n644_), .A2(new_n706_), .A3(new_n652_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n265_), .A2(G29gat), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT112), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n708_), .B2(new_n710_), .ZN(G1328gat));
  NAND3_X1  g510(.A1(new_n695_), .A2(new_n703_), .A3(new_n405_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G36gat), .ZN(new_n713_));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n707_), .A2(new_n714_), .A3(new_n405_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT45), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n713_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n713_), .A2(new_n716_), .A3(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  INV_X1    g520(.A(new_n455_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n695_), .A2(new_n703_), .A3(G43gat), .A4(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(G43gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n708_), .B2(new_n455_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n707_), .B2(new_n305_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n695_), .A2(new_n305_), .A3(new_n703_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G50gat), .ZN(G1331gat));
  INV_X1    g529(.A(new_n550_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(new_n584_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n467_), .A2(new_n732_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n733_), .A2(new_n639_), .A3(new_n653_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(G57gat), .A3(new_n264_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n643_), .B2(new_n733_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n640_), .A2(KEYINPUT113), .A3(new_n467_), .A4(new_n732_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n264_), .A3(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740_));
  INV_X1    g539(.A(G57gat), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n739_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n735_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT115), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n746_), .B(new_n735_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1332gat));
  NAND2_X1  g547(.A1(new_n734_), .A2(new_n405_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G64gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT48), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n737_), .A2(new_n738_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n405_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n753_), .A2(G64gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n752_), .B2(new_n754_), .ZN(G1333gat));
  INV_X1    g554(.A(G71gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n734_), .B2(new_n722_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT49), .Z(new_n758_));
  INV_X1    g557(.A(new_n752_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(new_n756_), .A3(new_n722_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1334gat));
  INV_X1    g560(.A(G78gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n734_), .B2(new_n305_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT50), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n759_), .A2(new_n762_), .A3(new_n305_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1335gat));
  NOR3_X1   g565(.A1(new_n733_), .A2(new_n706_), .A3(new_n652_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G85gat), .B1(new_n767_), .B2(new_n264_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT116), .B1(new_n701_), .B2(new_n702_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n693_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n731_), .A2(new_n706_), .A3(new_n584_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NOR4_X1   g574(.A1(new_n770_), .A2(new_n773_), .A3(new_n265_), .A4(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n768_), .B1(new_n776_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g576(.A(G92gat), .B1(new_n767_), .B2(new_n405_), .ZN(new_n778_));
  NOR4_X1   g577(.A1(new_n770_), .A2(new_n773_), .A3(new_n382_), .A4(new_n775_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n405_), .ZN(G1337gat));
  NAND4_X1  g579(.A1(new_n769_), .A2(new_n772_), .A3(new_n722_), .A4(new_n774_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G99gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n767_), .A2(new_n482_), .A3(new_n722_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT51), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n782_), .A2(new_n786_), .A3(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n767_), .A2(new_n473_), .A3(new_n305_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n305_), .B(new_n774_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(G106gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(G106gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n789_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  NAND4_X1  g597(.A1(new_n684_), .A2(new_n731_), .A3(new_n706_), .A4(new_n585_), .ZN(new_n799_));
  XOR2_X1   g598(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT118), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n639_), .B(new_n584_), .C1(new_n683_), .C2(new_n624_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  INV_X1    g602(.A(new_n800_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n731_), .A4(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n799_), .A2(new_n800_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n801_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n531_), .A2(new_n470_), .A3(new_n532_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n533_), .B1(KEYINPUT55), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n811_), .B(new_n470_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n538_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT56), .B(new_n538_), .C1(new_n810_), .C2(new_n812_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n813_), .A2(KEYINPUT121), .A3(new_n814_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n565_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n572_), .A2(new_n567_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n581_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n583_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n538_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n534_), .A2(new_n824_), .A3(new_n544_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n819_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n808_), .B1(new_n818_), .B2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(KEYINPUT58), .A3(new_n826_), .A4(new_n819_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n626_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n823_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n823_), .B(KEYINPUT119), .C1(new_n545_), .C2(new_n546_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n584_), .A2(new_n825_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT57), .B(new_n652_), .C1(new_n836_), .C2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n652_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n831_), .A2(new_n839_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n639_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n807_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n405_), .A2(new_n265_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n846_), .A2(new_n457_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G113gat), .B1(new_n849_), .B2(new_n584_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n831_), .A2(KEYINPUT123), .A3(new_n842_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n839_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT123), .B1(new_n831_), .B2(new_n842_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n639_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n807_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n847_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n848_), .A2(KEYINPUT59), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n584_), .A2(G113gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT124), .Z(new_n861_));
  AOI21_X1  g660(.A(new_n850_), .B1(new_n859_), .B2(new_n861_), .ZN(G1340gat));
  NAND3_X1  g661(.A1(new_n857_), .A2(new_n550_), .A3(new_n858_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G120gat), .ZN(new_n864_));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n731_), .B2(KEYINPUT60), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n849_), .B(new_n866_), .C1(KEYINPUT60), .C2(new_n865_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(G1341gat));
  NAND4_X1  g667(.A1(new_n857_), .A2(G127gat), .A3(new_n706_), .A4(new_n858_), .ZN(new_n869_));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n848_), .B2(new_n639_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1342gat));
  NAND4_X1  g671(.A1(new_n857_), .A2(G134gat), .A3(new_n626_), .A4(new_n858_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n233_), .B1(new_n848_), .B2(new_n652_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1343gat));
  AOI211_X1 g674(.A(new_n429_), .B(new_n722_), .C1(new_n807_), .C2(new_n844_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n584_), .A3(new_n846_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n550_), .A3(new_n846_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g679(.A1(new_n876_), .A2(new_n706_), .A3(new_n846_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  AND2_X1   g682(.A1(new_n876_), .A2(new_n846_), .ZN(new_n884_));
  INV_X1    g683(.A(G162gat), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n698_), .A2(new_n699_), .A3(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n876_), .A2(new_n653_), .A3(new_n846_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n884_), .A2(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1347gat));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n753_), .A2(new_n264_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n457_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n585_), .B(new_n892_), .C1(new_n854_), .C2(new_n807_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n889_), .B(new_n890_), .C1(new_n893_), .C2(new_n317_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n892_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n855_), .A2(new_n584_), .A3(new_n895_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n896_), .A2(new_n367_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n889_), .A2(new_n890_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n896_), .A2(G169gat), .A3(new_n898_), .A4(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n894_), .A2(new_n897_), .A3(new_n900_), .ZN(G1348gat));
  NAND3_X1  g700(.A1(new_n845_), .A2(new_n550_), .A3(new_n895_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G176gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n855_), .A2(new_n895_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n731_), .A2(G176gat), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n903_), .B1(new_n904_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT126), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n903_), .B(new_n909_), .C1(new_n904_), .C2(new_n906_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1349gat));
  NOR3_X1   g710(.A1(new_n904_), .A2(new_n639_), .A3(new_n307_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n845_), .A2(new_n706_), .A3(new_n895_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n322_), .B2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n904_), .B2(new_n684_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n653_), .A2(new_n359_), .A3(new_n309_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n904_), .B2(new_n916_), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n876_), .A2(new_n584_), .A3(new_n891_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g718(.A1(new_n876_), .A2(new_n550_), .A3(new_n891_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n876_), .A2(new_n891_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n639_), .ZN(new_n924_));
  XOR2_X1   g723(.A(KEYINPUT63), .B(G211gat), .Z(new_n925_));
  NAND4_X1  g724(.A1(new_n876_), .A2(new_n706_), .A3(new_n891_), .A4(new_n925_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1354gat));
  INV_X1    g726(.A(G218gat), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n923_), .A2(new_n928_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n876_), .A2(new_n653_), .A3(new_n891_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n929_), .A2(new_n626_), .B1(new_n928_), .B2(new_n930_), .ZN(G1355gat));
endmodule


