//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT74), .ZN(new_n203_));
  XOR2_X1   g002(.A(G134gat), .B(G162gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT36), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G232gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT34), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT35), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT6), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT6), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n218_), .A2(new_n220_), .A3(KEYINPUT66), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT68), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT67), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n230_), .B1(KEYINPUT68), .B2(new_n226_), .ZN(new_n231_));
  OAI22_X1  g030(.A1(KEYINPUT67), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n229_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n216_), .B1(new_n225_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n214_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(new_n233_), .B2(new_n221_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n215_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT67), .B1(new_n239_), .B2(KEYINPUT7), .ZN(new_n240_));
  INV_X1    g039(.A(G99gat), .ZN(new_n241_));
  INV_X1    g040(.A(G106gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n230_), .A2(new_n226_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n245_), .A2(new_n229_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT69), .B1(new_n246_), .B2(new_n235_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n234_), .B1(new_n238_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT10), .B(G99gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n225_), .B1(G106gat), .B2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n213_), .B1(new_n212_), .B2(KEYINPUT9), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT9), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n211_), .A2(KEYINPUT64), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT64), .B1(new_n211_), .B2(new_n252_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n251_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT65), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n255_), .A2(KEYINPUT65), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n250_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n248_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G43gat), .B(G50gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G29gat), .B(G36gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT73), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n262_), .A2(KEYINPUT73), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n261_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n265_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(new_n263_), .A3(new_n260_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n210_), .B1(new_n259_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n209_), .A2(KEYINPUT35), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT72), .Z(new_n272_));
  NOR2_X1   g071(.A1(new_n231_), .A2(new_n232_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n240_), .A2(new_n243_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n221_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(new_n237_), .A3(new_n214_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n247_), .A2(new_n276_), .A3(KEYINPUT8), .ZN(new_n277_));
  INV_X1    g076(.A(new_n234_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT71), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n281_), .A3(new_n278_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n258_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT15), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n269_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n266_), .A2(new_n268_), .A3(KEYINPUT15), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n270_), .B(new_n272_), .C1(new_n283_), .C2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n258_), .ZN(new_n290_));
  AOI211_X1 g089(.A(KEYINPUT71), .B(new_n234_), .C1(new_n238_), .C2(new_n247_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n281_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n287_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n272_), .B1(new_n295_), .B2(new_n270_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n206_), .A2(KEYINPUT36), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n289_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n270_), .B1(new_n283_), .B2(new_n287_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n272_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n297_), .B1(new_n302_), .B2(new_n288_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n207_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n297_), .A3(new_n288_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT37), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n298_), .B1(new_n289_), .B2(new_n296_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n305_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n311_), .A2(KEYINPUT37), .A3(new_n307_), .A4(new_n207_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G127gat), .B(G155gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT16), .ZN(new_n315_));
  XOR2_X1   g114(.A(G183gat), .B(G211gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT17), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G57gat), .B(G64gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G71gat), .B(G78gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(KEYINPUT11), .ZN(new_n322_));
  XOR2_X1   g121(.A(G71gat), .B(G78gat), .Z(new_n323_));
  INV_X1    g122(.A(G64gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G57gat), .ZN(new_n325_));
  INV_X1    g124(.A(G57gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G64gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n327_), .A3(KEYINPUT11), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n320_), .A2(KEYINPUT11), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n322_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT77), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G15gat), .B(G22gat), .ZN(new_n335_));
  INV_X1    g134(.A(G1gat), .ZN(new_n336_));
  INV_X1    g135(.A(G8gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT14), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G1gat), .B(G8gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G231gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n319_), .B1(new_n334_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n343_), .B2(new_n334_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n343_), .A2(new_n331_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n317_), .A2(new_n318_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n331_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n349_), .A2(KEYINPUT76), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(KEYINPUT76), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n313_), .A2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n354_), .B(KEYINPUT78), .Z(new_n355_));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT19), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G169gat), .ZN(new_n358_));
  INV_X1    g157(.A(G176gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT83), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT96), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(G183gat), .A3(G190gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(G183gat), .B2(G190gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n370_), .A2(KEYINPUT84), .ZN(new_n371_));
  INV_X1    g170(.A(G183gat), .ZN(new_n372_));
  INV_X1    g171(.A(G190gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT23), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n369_), .B1(new_n371_), .B2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT25), .B(G183gat), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n381_), .A2(KEYINPUT95), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT26), .B(G190gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(KEYINPUT95), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n374_), .A2(new_n369_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n361_), .B2(new_n391_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n367_), .A2(new_n380_), .B1(new_n385_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G211gat), .B(G218gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT21), .ZN(new_n396_));
  INV_X1    g195(.A(G197gat), .ZN(new_n397_));
  INV_X1    g196(.A(G204gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT93), .B(G197gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(new_n398_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n398_), .A2(G197gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT94), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n400_), .A2(G204gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT21), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT21), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n395_), .B1(new_n401_), .B2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n402_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT20), .B1(new_n393_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT85), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n377_), .A2(new_n411_), .A3(new_n388_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n369_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n370_), .A2(KEYINPUT84), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n374_), .A2(new_n375_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT85), .B1(new_n416_), .B2(new_n387_), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n362_), .A2(new_n391_), .B1(new_n383_), .B2(new_n381_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n412_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n386_), .A2(new_n379_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT22), .ZN(new_n421_));
  OAI21_X1  g220(.A(G169gat), .B1(new_n421_), .B2(KEYINPUT86), .ZN(new_n422_));
  INV_X1    g221(.A(G169gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT22), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n422_), .B(new_n359_), .C1(KEYINPUT86), .C2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n420_), .A2(new_n425_), .A3(new_n362_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n419_), .A2(new_n409_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n357_), .B1(new_n410_), .B2(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G8gat), .B(G36gat), .Z(new_n430_));
  XNOR2_X1  g229(.A(G64gat), .B(G92gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n393_), .B2(new_n409_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n419_), .A2(new_n426_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n409_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n357_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n429_), .A2(new_n434_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT27), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n434_), .B(KEYINPUT102), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n366_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n380_), .A2(new_n446_), .A3(new_n364_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n392_), .A2(new_n385_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n435_), .B1(new_n449_), .B2(new_n438_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(new_n440_), .A3(new_n427_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT20), .B1(new_n449_), .B2(new_n438_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n409_), .B1(new_n419_), .B2(new_n426_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n357_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n445_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT103), .B1(new_n443_), .B2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(G155gat), .A2(G162gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT1), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n457_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT90), .B1(G141gat), .B2(G148gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(KEYINPUT90), .A2(G141gat), .A3(G148gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n461_), .B(new_n462_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  OR3_X1    g265(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT2), .ZN(new_n468_));
  INV_X1    g267(.A(G141gat), .ZN(new_n469_));
  INV_X1    g268(.A(G148gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n467_), .A2(new_n471_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n459_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n466_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT92), .B1(new_n476_), .B2(KEYINPUT29), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n438_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G228gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(G78gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(G106gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n478_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT28), .B1(new_n476_), .B2(KEYINPUT29), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n476_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT91), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n487_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n485_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G22gat), .B(G50gat), .Z(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n488_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n484_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(new_n494_), .A3(new_n483_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n434_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n452_), .A2(new_n357_), .A3(new_n453_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n440_), .B1(new_n450_), .B2(new_n427_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n442_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT27), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n451_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n440_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n444_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT103), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT27), .A4(new_n442_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n456_), .A2(new_n500_), .A3(new_n507_), .A4(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G227gat), .A2(G233gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n514_), .B(G71gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(new_n241_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n437_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G15gat), .B(G43gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT87), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT30), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n437_), .A2(new_n516_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n518_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n522_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n523_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n521_), .B1(new_n529_), .B2(new_n517_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT89), .B1(new_n530_), .B2(new_n524_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G113gat), .B(G120gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G127gat), .B(G134gat), .Z(new_n534_));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G127gat), .B(G134gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT88), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n533_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n535_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(KEYINPUT88), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(new_n541_), .A3(new_n532_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT31), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n528_), .A2(new_n531_), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(KEYINPUT98), .A3(new_n476_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n539_), .A2(new_n466_), .A3(new_n475_), .A4(new_n542_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(KEYINPUT4), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT4), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n543_), .A2(KEYINPUT98), .A3(new_n549_), .A4(new_n476_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G225gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G1gat), .B(G29gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(G85gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT0), .B(G57gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n543_), .A2(new_n476_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n547_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n552_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n554_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n558_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n552_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n561_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n562_), .A2(KEYINPUT101), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT101), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n554_), .A2(new_n568_), .A3(new_n558_), .A4(new_n561_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n544_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT89), .B(new_n571_), .C1(new_n530_), .C2(new_n524_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n545_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n513_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n434_), .A2(KEYINPUT32), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n429_), .A2(new_n441_), .A3(new_n575_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n567_), .A2(new_n569_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(KEYINPUT33), .B(new_n563_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT33), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n566_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n558_), .B1(new_n560_), .B2(new_n552_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT100), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT100), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n587_), .B(new_n558_), .C1(new_n560_), .C2(new_n552_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n586_), .B(new_n588_), .C1(new_n553_), .C2(new_n551_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n584_), .A2(new_n504_), .A3(new_n442_), .A4(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n579_), .B1(new_n582_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n500_), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n569_), .A2(new_n567_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n593_), .A2(new_n456_), .A3(new_n507_), .A4(new_n512_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n545_), .A2(new_n572_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n574_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n248_), .A2(new_n333_), .A3(new_n258_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n333_), .B1(new_n248_), .B2(new_n258_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n331_), .A2(new_n600_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n293_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G230gat), .A2(G233gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n601_), .ZN(new_n608_));
  OAI211_X1 g407(.A(G230gat), .B(G233gat), .C1(new_n608_), .C2(new_n599_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT5), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n607_), .A2(new_n609_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n598_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(KEYINPUT13), .A3(new_n615_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n341_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n269_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n341_), .A2(new_n268_), .A3(new_n266_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(KEYINPUT79), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT79), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n341_), .A2(new_n268_), .A3(new_n266_), .A4(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n269_), .B2(new_n622_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n631_), .B1(new_n287_), .B2(new_n622_), .ZN(new_n632_));
  XOR2_X1   g431(.A(G113gat), .B(G141gat), .Z(new_n633_));
  XOR2_X1   g432(.A(G169gat), .B(G197gat), .Z(new_n634_));
  XOR2_X1   g433(.A(new_n633_), .B(new_n634_), .Z(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(new_n632_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT81), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT81), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n630_), .A2(new_n632_), .A3(new_n638_), .A4(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n635_), .B(KEYINPUT80), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT82), .B1(new_n640_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT82), .ZN(new_n645_));
  AOI211_X1 g444(.A(new_n645_), .B(new_n642_), .C1(new_n637_), .C2(new_n639_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n597_), .A2(new_n621_), .A3(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n355_), .A2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n570_), .B(KEYINPUT104), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n336_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n621_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n640_), .A2(new_n643_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n353_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n597_), .A2(new_n304_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(new_n657_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n570_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n651_), .A2(new_n652_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n653_), .A2(new_n662_), .A3(new_n663_), .ZN(G1324gat));
  NAND3_X1  g463(.A1(new_n456_), .A2(new_n507_), .A3(new_n512_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n649_), .A2(new_n337_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  INV_X1    g466(.A(new_n661_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n665_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n669_), .B2(G8gat), .ZN(new_n670_));
  AOI211_X1 g469(.A(KEYINPUT39), .B(new_n337_), .C1(new_n668_), .C2(new_n665_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g472(.A(G15gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n596_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n649_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n668_), .A2(new_n675_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n677_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT41), .B1(new_n677_), .B2(G15gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n500_), .A2(G22gat), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT106), .Z(new_n682_));
  NAND2_X1  g481(.A1(new_n649_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G22gat), .B1(new_n661_), .B2(new_n500_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(KEYINPUT42), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(KEYINPUT42), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(G1327gat));
  INV_X1    g486(.A(new_n304_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(new_n353_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n648_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n570_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G29gat), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n655_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n621_), .A2(new_n353_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n456_), .A2(new_n507_), .A3(new_n512_), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n697_), .A2(new_n593_), .B1(new_n591_), .B2(new_n500_), .ZN(new_n698_));
  OAI22_X1  g497(.A1(new_n698_), .A2(new_n675_), .B1(new_n513_), .B2(new_n573_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n313_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n597_), .A2(KEYINPUT43), .A3(new_n313_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n695_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT107), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  INV_X1    g504(.A(new_n695_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n699_), .A2(new_n700_), .A3(new_n696_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n597_), .B2(new_n313_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n706_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n704_), .A2(new_n705_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(KEYINPUT44), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n650_), .A2(G29gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n693_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  NAND3_X1  g515(.A1(new_n712_), .A2(new_n665_), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n665_), .B(KEYINPUT108), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n690_), .A2(G36gat), .A3(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(KEYINPUT46), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n718_), .B(new_n723_), .C1(new_n725_), .C2(KEYINPUT46), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1329gat));
  INV_X1    g528(.A(G43gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n730_), .B1(new_n690_), .B2(new_n596_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n675_), .A2(G43gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n709_), .B2(KEYINPUT44), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n712_), .B2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT107), .B(new_n706_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n732_), .B(new_n734_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n731_), .B1(new_n735_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT47), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n742_), .B(new_n731_), .C1(new_n735_), .C2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1330gat));
  OR3_X1    g543(.A1(new_n690_), .A2(G50gat), .A3(new_n500_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n500_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n712_), .A2(new_n746_), .A3(new_n713_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(KEYINPUT112), .ZN(new_n748_));
  OAI21_X1  g547(.A(G50gat), .B1(new_n747_), .B2(KEYINPUT112), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1331gat));
  NOR3_X1   g549(.A1(new_n644_), .A2(new_n646_), .A3(new_n352_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n659_), .A2(new_n621_), .A3(new_n751_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n752_), .A2(new_n326_), .A3(new_n570_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n597_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n355_), .A2(new_n754_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n755_), .A2(KEYINPUT113), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(KEYINPUT113), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n650_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n753_), .B1(new_n758_), .B2(new_n326_), .ZN(G1332gat));
  OAI21_X1  g558(.A(G64gat), .B1(new_n752_), .B2(new_n720_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT48), .ZN(new_n761_));
  INV_X1    g560(.A(new_n755_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n324_), .A3(new_n719_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1333gat));
  OAI21_X1  g563(.A(G71gat), .B1(new_n752_), .B2(new_n596_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT49), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n596_), .A2(G71gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n755_), .B2(new_n767_), .ZN(G1334gat));
  OAI21_X1  g567(.A(G78gat), .B1(new_n752_), .B2(new_n500_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n770_));
  XNOR2_X1  g569(.A(new_n769_), .B(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n762_), .A2(new_n480_), .A3(new_n746_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1335gat));
  NAND2_X1  g572(.A1(new_n754_), .A2(new_n689_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(G85gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n650_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n621_), .A2(new_n352_), .A3(new_n694_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(new_n692_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n780_), .B2(new_n776_), .ZN(G1336gat));
  INV_X1    g580(.A(G92gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n775_), .A2(new_n782_), .A3(new_n665_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n779_), .A2(new_n719_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n782_), .ZN(G1337gat));
  AOI21_X1  g584(.A(new_n241_), .B1(new_n779_), .B2(new_n675_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n774_), .A2(new_n249_), .A3(new_n596_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g588(.A1(new_n779_), .A2(KEYINPUT116), .A3(new_n746_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n790_), .A2(G106gat), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n779_), .A2(new_n746_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(KEYINPUT52), .A3(new_n794_), .ZN(new_n795_));
  AND4_X1   g594(.A1(new_n242_), .A2(new_n754_), .A3(new_n746_), .A4(new_n689_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT115), .Z(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(new_n791_), .B2(new_n794_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT53), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n799_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n795_), .A4(new_n797_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n803_), .ZN(G1339gat));
  AND3_X1   g603(.A1(new_n751_), .A2(new_n620_), .A3(new_n618_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n313_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n313_), .B(new_n805_), .C1(KEYINPUT117), .C2(KEYINPUT54), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n808_), .A2(new_n809_), .B1(KEYINPUT117), .B2(KEYINPUT54), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n655_), .A2(new_n615_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n606_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n607_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n602_), .A2(new_n605_), .A3(KEYINPUT55), .A4(new_n606_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n613_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(KEYINPUT56), .A3(new_n613_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n811_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n625_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n635_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n287_), .A2(new_n622_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n623_), .A2(new_n629_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n823_), .B(new_n824_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n640_), .A2(new_n822_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n822_), .B1(new_n640_), .B2(new_n827_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n619_), .B2(new_n615_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n688_), .B1(new_n821_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT57), .B(new_n688_), .C1(new_n821_), .C2(new_n831_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n615_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n816_), .B2(new_n613_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n818_), .B(new_n614_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n313_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n837_), .B(KEYINPUT58), .C1(new_n838_), .C2(new_n839_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n834_), .A2(new_n835_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n810_), .B1(new_n845_), .B2(new_n352_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n513_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n650_), .A2(new_n675_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(KEYINPUT120), .ZN(new_n850_));
  OR3_X1    g649(.A1(new_n846_), .A2(new_n848_), .A3(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n849_), .A2(KEYINPUT120), .ZN(new_n852_));
  OAI22_X1  g651(.A1(new_n846_), .A2(new_n848_), .B1(new_n852_), .B2(new_n850_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G113gat), .B1(new_n854_), .B2(new_n647_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n848_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n832_), .A2(new_n833_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n353_), .B1(new_n859_), .B2(new_n835_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT119), .B(new_n858_), .C1(new_n860_), .C2(new_n810_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n694_), .A2(G113gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n857_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n855_), .A2(new_n863_), .ZN(G1340gat));
  OAI21_X1  g663(.A(G120gat), .B1(new_n854_), .B2(new_n654_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT60), .ZN(new_n866_));
  AOI21_X1  g665(.A(G120gat), .B1(new_n621_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(G120gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(KEYINPUT121), .B2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(KEYINPUT121), .B2(new_n867_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n857_), .A2(new_n861_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n865_), .A2(new_n871_), .ZN(G1341gat));
  OAI21_X1  g671(.A(G127gat), .B1(new_n854_), .B2(new_n352_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n352_), .A2(G127gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n857_), .A2(new_n861_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1342gat));
  AND4_X1   g675(.A1(G134gat), .A2(new_n851_), .A3(new_n700_), .A4(new_n853_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n857_), .A2(new_n304_), .A3(new_n861_), .ZN(new_n878_));
  INV_X1    g677(.A(G134gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT122), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n878_), .A2(new_n882_), .A3(new_n879_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n877_), .B1(new_n881_), .B2(new_n883_), .ZN(G1343gat));
  INV_X1    g683(.A(new_n846_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n675_), .A2(new_n500_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n885_), .A2(new_n650_), .A3(new_n720_), .A4(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n694_), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT123), .B(G141gat), .Z(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n887_), .A2(new_n654_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n470_), .ZN(G1345gat));
  NOR2_X1   g691(.A1(new_n887_), .A2(new_n352_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n893_), .B(new_n895_), .ZN(G1346gat));
  OAI21_X1  g695(.A(G162gat), .B1(new_n887_), .B2(new_n313_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n688_), .A2(G162gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n887_), .B2(new_n898_), .ZN(G1347gat));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n650_), .A2(new_n596_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n719_), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT124), .Z(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n500_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n846_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n694_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n900_), .B1(new_n907_), .B2(new_n423_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n358_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT62), .B(G169gat), .C1(new_n906_), .C2(new_n694_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n909_), .A3(new_n910_), .ZN(G1348gat));
  NAND2_X1  g710(.A1(new_n905_), .A2(new_n621_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g712(.A1(new_n905_), .A2(new_n353_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n382_), .A2(new_n384_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n914_), .A2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G183gat), .B1(new_n905_), .B2(new_n353_), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT125), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n914_), .A2(new_n372_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n920_), .B(new_n921_), .C1(new_n916_), .C2(new_n914_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n919_), .A2(new_n922_), .ZN(G1350gat));
  OAI21_X1  g722(.A(G190gat), .B1(new_n906_), .B2(new_n313_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n905_), .A2(new_n304_), .A3(new_n383_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1351gat));
  NAND2_X1  g725(.A1(new_n596_), .A2(new_n593_), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT126), .Z(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n720_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n885_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n694_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(new_n397_), .ZN(G1352gat));
  NOR2_X1   g731(.A1(new_n930_), .A2(new_n654_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n398_), .ZN(G1353gat));
  NOR2_X1   g733(.A1(new_n930_), .A2(new_n352_), .ZN(new_n935_));
  OR2_X1    g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT63), .B(G211gat), .Z(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n935_), .B2(new_n938_), .ZN(G1354gat));
  INV_X1    g738(.A(G218gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n930_), .A2(new_n940_), .A3(new_n313_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n930_), .A2(KEYINPUT127), .A3(new_n688_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(G218gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(KEYINPUT127), .B1(new_n930_), .B2(new_n688_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n941_), .B1(new_n943_), .B2(new_n944_), .ZN(G1355gat));
endmodule


