//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n208_), .B(new_n209_), .C1(new_n212_), .C2(KEYINPUT24), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(G169gat), .B2(G176gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT77), .ZN(new_n217_));
  INV_X1    g016(.A(G190gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n217_), .B1(new_n218_), .B2(KEYINPUT26), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n219_), .B(new_n220_), .C1(new_n221_), .C2(new_n217_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(G169gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n208_), .B(new_n209_), .C1(G183gat), .C2(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT21), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(KEYINPUT21), .A3(new_n230_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n234_), .A2(new_n235_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n228_), .A2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n213_), .A2(KEYINPUT85), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n213_), .A2(KEYINPUT85), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n215_), .B1(new_n221_), .B2(new_n220_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n236_), .A2(new_n237_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n227_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT87), .ZN(new_n246_));
  OAI211_X1 g045(.A(KEYINPUT20), .B(new_n239_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n245_), .A2(new_n246_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n205_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(new_n227_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n238_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT86), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n250_), .A2(KEYINPUT86), .A3(new_n238_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT20), .ZN(new_n255_));
  INV_X1    g054(.A(new_n228_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(new_n244_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n253_), .A2(new_n204_), .A3(new_n254_), .A4(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n249_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT89), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G8gat), .B(G36gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G64gat), .B(G92gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n263_), .B(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n259_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n263_), .B(new_n264_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n249_), .A2(new_n258_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT27), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT99), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT99), .ZN(new_n274_));
  INV_X1    g073(.A(new_n269_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n268_), .B1(new_n249_), .B2(new_n258_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n274_), .B(new_n271_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G113gat), .B(G120gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G127gat), .B(G134gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT78), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n281_), .A2(KEYINPUT78), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n280_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n281_), .A2(KEYINPUT78), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(new_n282_), .A3(new_n279_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G71gat), .B(G99gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(G43gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n228_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G227gat), .A2(G233gat), .ZN(new_n294_));
  INV_X1    g093(.A(G15gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT30), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n297_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n290_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT80), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n301_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n298_), .A2(new_n299_), .A3(new_n290_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT81), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(KEYINPUT81), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n302_), .A2(new_n303_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G1gat), .B(G29gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT95), .B(G85gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT0), .B(G57gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT93), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT1), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT82), .ZN(new_n317_));
  OR2_X1    g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(new_n319_), .A3(KEYINPUT1), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(G155gat), .A3(G162gat), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n317_), .A2(new_n318_), .A3(new_n320_), .A4(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  INV_X1    g123(.A(G141gat), .ZN(new_n325_));
  INV_X1    g124(.A(G148gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n323_), .A2(new_n324_), .A3(new_n327_), .ZN(new_n328_));
  OR3_X1    g127(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n318_), .A2(new_n315_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT83), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT83), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n318_), .A2(new_n337_), .A3(new_n315_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n328_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(KEYINPUT94), .B(KEYINPUT4), .Z(new_n341_));
  NAND3_X1  g140(.A1(new_n288_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n328_), .A2(new_n339_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT92), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n287_), .A4(new_n285_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT92), .B1(new_n288_), .B2(new_n340_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n288_), .A2(new_n340_), .A3(KEYINPUT91), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT91), .B1(new_n288_), .B2(new_n340_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n345_), .B(new_n346_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n314_), .B(new_n342_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n347_), .A2(new_n348_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n314_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n346_), .A4(new_n345_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n312_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(new_n354_), .A3(new_n312_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n307_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n253_), .A2(new_n205_), .A3(new_n254_), .A4(new_n257_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n360_), .A2(KEYINPUT98), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n362_));
  NAND3_X1  g161(.A1(new_n245_), .A2(new_n239_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n204_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(KEYINPUT98), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n268_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n276_), .A2(new_n271_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT84), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n343_), .B2(new_n372_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n340_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G22gat), .B(G50gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n373_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n343_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT28), .B1(new_n340_), .B2(KEYINPUT29), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n370_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n244_), .B1(new_n340_), .B2(KEYINPUT29), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383_));
  INV_X1    g182(.A(G78gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G106gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n382_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n376_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n378_), .A2(new_n379_), .A3(new_n375_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(KEYINPUT84), .A3(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n381_), .A2(new_n388_), .A3(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n387_), .B(new_n370_), .C1(new_n377_), .C2(new_n380_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AND4_X1   g193(.A1(new_n278_), .A2(new_n359_), .A3(new_n369_), .A4(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n267_), .A2(KEYINPUT90), .A3(new_n269_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n349_), .A2(new_n353_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(new_n312_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n353_), .B(new_n342_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n357_), .A2(new_n400_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n357_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT33), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n366_), .A2(KEYINPUT32), .A3(new_n266_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT96), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n266_), .A2(KEYINPUT32), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n259_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n259_), .B2(new_n410_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n358_), .A2(new_n408_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n407_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n394_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n405_), .A2(new_n394_), .A3(new_n355_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n274_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n277_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n417_), .B(new_n369_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT100), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n278_), .A2(KEYINPUT100), .A3(new_n369_), .A4(new_n417_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n416_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n395_), .B1(new_n424_), .B2(new_n307_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT70), .ZN(new_n426_));
  XOR2_X1   g225(.A(G29gat), .B(G36gat), .Z(new_n427_));
  XOR2_X1   g226(.A(G43gat), .B(G50gat), .Z(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G29gat), .B(G36gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G43gat), .B(G50gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(KEYINPUT15), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT15), .B1(new_n429_), .B2(new_n432_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n437_));
  INV_X1    g236(.A(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(G85gat), .A2(G92gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(KEYINPUT9), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G99gat), .A2(G106gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT6), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n442_), .A2(KEYINPUT9), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n440_), .A2(new_n443_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n441_), .A2(new_n442_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI211_X1 g254(.A(KEYINPUT8), .B(new_n451_), .C1(new_n455_), .C2(new_n448_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT8), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT7), .ZN(new_n458_));
  INV_X1    g257(.A(G99gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n438_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n448_), .A2(new_n452_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n451_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n457_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n450_), .B1(new_n456_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n436_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G232gat), .A2(G233gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT34), .Z(new_n467_));
  XOR2_X1   g266(.A(KEYINPUT66), .B(KEYINPUT35), .Z(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n469_), .B(KEYINPUT69), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n468_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n429_), .A2(new_n432_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n464_), .B2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n426_), .B1(new_n471_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n450_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n445_), .A2(new_n447_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n460_), .A2(new_n452_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n462_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT8), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n461_), .A2(new_n457_), .A3(new_n462_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n477_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n483_), .A2(new_n473_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n484_), .A2(KEYINPUT70), .A3(new_n465_), .A4(new_n470_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n476_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT68), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n465_), .A2(KEYINPUT67), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT67), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n436_), .A2(new_n464_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n484_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n469_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n486_), .A2(new_n487_), .A3(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G190gat), .B(G218gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G134gat), .B(G162gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(KEYINPUT36), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n486_), .A2(new_n487_), .A3(new_n492_), .A4(new_n497_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n486_), .A2(new_n492_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(KEYINPUT36), .A3(new_n496_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n425_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G120gat), .B(G148gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT64), .B(KEYINPUT5), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G176gat), .B(G204gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G64gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G71gat), .B(G78gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT11), .ZN(new_n514_));
  INV_X1    g313(.A(new_n513_), .ZN(new_n515_));
  INV_X1    g314(.A(G64gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(G57gat), .ZN(new_n517_));
  INV_X1    g316(.A(G57gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(G64gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n519_), .A3(KEYINPUT11), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n512_), .A2(KEYINPUT11), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n514_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n450_), .B(new_n523_), .C1(new_n456_), .C2(new_n463_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G230gat), .A2(G233gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT12), .B1(new_n483_), .B2(new_n523_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n528_));
  INV_X1    g327(.A(new_n523_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n464_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n526_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n464_), .A2(new_n529_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n525_), .B1(new_n532_), .B2(new_n524_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n511_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n525_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(new_n483_), .B2(new_n523_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n483_), .A2(KEYINPUT12), .A3(new_n523_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n528_), .B1(new_n464_), .B2(new_n529_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n536_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n532_), .A2(new_n524_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n535_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n541_), .A3(new_n510_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT65), .B1(new_n534_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT13), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n534_), .A2(new_n542_), .A3(KEYINPUT65), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n534_), .A2(new_n542_), .A3(KEYINPUT65), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT13), .B1(new_n548_), .B2(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(G8gat), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n295_), .A2(KEYINPUT71), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT71), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(G15gat), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n554_), .A2(new_n556_), .A3(G22gat), .ZN(new_n557_));
  AOI21_X1  g356(.A(G22gat), .B1(new_n554_), .B2(new_n556_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n553_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G1gat), .B(G8gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n554_), .A2(new_n556_), .ZN(new_n562_));
  INV_X1    g361(.A(G22gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n554_), .A2(new_n556_), .A3(G22gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n560_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n553_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n561_), .A2(new_n568_), .A3(new_n473_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT76), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n567_), .B1(new_n566_), .B2(new_n553_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n553_), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n560_), .B(new_n576_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT15), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n473_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n433_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n578_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n561_), .A2(new_n568_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT75), .B1(new_n436_), .B2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n574_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n474_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n569_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(G229gat), .A3(G233gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G169gat), .B(G197gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n586_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n578_), .B(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n600_), .A2(new_n523_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n584_), .B(new_n599_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(new_n529_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT73), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT16), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT17), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n600_), .A2(new_n523_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT73), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n602_), .A2(new_n529_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n608_), .A2(KEYINPUT17), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n604_), .A2(new_n609_), .A3(new_n613_), .A4(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n609_), .B(KEYINPUT72), .Z(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n551_), .A2(new_n598_), .A3(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n505_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n202_), .B1(new_n620_), .B2(new_n358_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT102), .Z(new_n622_));
  NOR3_X1   g421(.A1(new_n425_), .A2(new_n598_), .A3(new_n551_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT37), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n501_), .A2(new_n624_), .A3(new_n503_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n618_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT74), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n623_), .A2(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n358_), .A2(KEYINPUT101), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n358_), .A2(KEYINPUT101), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n631_), .A2(new_n202_), .A3(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT38), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n622_), .A2(new_n636_), .ZN(G1324gat));
  NAND2_X1  g436(.A1(new_n278_), .A2(new_n369_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n631_), .A2(new_n552_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n620_), .A2(new_n638_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(G8gat), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n640_), .B2(G8gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(G1325gat));
  INV_X1    g445(.A(new_n307_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n295_), .B1(new_n620_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT41), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n631_), .A2(new_n295_), .A3(new_n647_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(new_n394_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n563_), .B1(new_n620_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n631_), .A2(new_n563_), .A3(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1327gat));
  NAND2_X1  g456(.A1(new_n424_), .A2(new_n307_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n395_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n551_), .A2(new_n598_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n504_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n628_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G29gat), .B1(new_n665_), .B2(new_n358_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n504_), .A2(KEYINPUT37), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n501_), .A2(new_n624_), .A3(new_n503_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n667_), .B1(new_n660_), .B2(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n425_), .A2(KEYINPUT43), .A3(new_n627_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n661_), .B(new_n618_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n660_), .A2(new_n667_), .A3(new_n670_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n425_), .B2(new_n627_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n678_), .A2(KEYINPUT44), .A3(new_n661_), .A4(new_n618_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n675_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n634_), .A2(G29gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n666_), .B1(new_n680_), .B2(new_n681_), .ZN(G1328gat));
  XNOR2_X1  g481(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n675_), .A2(new_n638_), .A3(new_n679_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  INV_X1    g484(.A(new_n638_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(G36gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT45), .B1(new_n664_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT45), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n623_), .A2(new_n690_), .A3(new_n663_), .A4(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n683_), .B1(new_n685_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n692_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n683_), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n694_), .B(new_n695_), .C1(new_n684_), .C2(G36gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1329gat));
  NAND4_X1  g496(.A1(new_n675_), .A2(G43gat), .A3(new_n647_), .A4(new_n679_), .ZN(new_n698_));
  INV_X1    g497(.A(G43gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n699_), .B1(new_n664_), .B2(new_n307_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g501(.A1(new_n664_), .A2(G50gat), .A3(new_n394_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n680_), .B2(new_n652_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n675_), .A2(new_n704_), .A3(new_n652_), .A4(new_n679_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G50gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n705_), .B2(new_n707_), .ZN(G1331gat));
  NOR2_X1   g507(.A1(new_n550_), .A2(new_n597_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n425_), .A2(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n630_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G57gat), .B1(new_n712_), .B2(new_n634_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n615_), .A2(new_n595_), .A3(new_n596_), .A4(new_n617_), .ZN(new_n714_));
  NOR4_X1   g513(.A1(new_n425_), .A2(new_n504_), .A3(new_n550_), .A4(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n358_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT107), .B(G57gat), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n713_), .B1(new_n715_), .B2(new_n718_), .ZN(G1332gat));
  AOI21_X1  g518(.A(new_n516_), .B1(new_n715_), .B2(new_n638_), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n712_), .A2(new_n516_), .A3(new_n638_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1333gat));
  INV_X1    g523(.A(G71gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n715_), .B2(new_n647_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n712_), .A2(new_n725_), .A3(new_n647_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1334gat));
  AOI21_X1  g529(.A(new_n384_), .B1(new_n715_), .B2(new_n652_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT50), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n712_), .A2(new_n384_), .A3(new_n652_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1335gat));
  AOI211_X1 g533(.A(new_n628_), .B(new_n710_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n358_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G85gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n711_), .A2(new_n663_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n634_), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n739_), .A2(G85gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n738_), .B2(new_n740_), .ZN(G1336gat));
  INV_X1    g540(.A(G92gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n742_), .B1(new_n738_), .B2(new_n686_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT110), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n638_), .A2(G92gat), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT111), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n735_), .B2(new_n746_), .ZN(G1337gat));
  NAND3_X1  g546(.A1(new_n647_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n738_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n735_), .A2(new_n647_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G99gat), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT51), .Z(G1338gat));
  NAND4_X1  g551(.A1(new_n711_), .A2(new_n438_), .A3(new_n652_), .A4(new_n663_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n678_), .A2(new_n652_), .A3(new_n618_), .A4(new_n709_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n755_), .A3(G106gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G106gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n753_), .B(new_n759_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1339gat));
  NOR4_X1   g562(.A1(new_n739_), .A2(new_n307_), .A3(new_n638_), .A4(new_n652_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT119), .ZN(new_n765_));
  INV_X1    g564(.A(new_n524_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n768_));
  OAI22_X1  g567(.A1(new_n525_), .A2(new_n767_), .B1(new_n531_), .B2(new_n768_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n531_), .A2(KEYINPUT55), .ZN(new_n770_));
  OAI211_X1 g569(.A(KEYINPUT56), .B(new_n511_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n768_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n539_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n531_), .A2(KEYINPUT55), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n775_), .B(new_n776_), .C1(new_n525_), .C2(new_n767_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n511_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n773_), .A2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n511_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(KEYINPUT114), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n542_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n779_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n473_), .B1(new_n561_), .B2(new_n568_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n572_), .B1(new_n570_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n594_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n569_), .A2(new_n573_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n582_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n436_), .A2(KEYINPUT75), .A3(new_n584_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT115), .B1(new_n789_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n790_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n593_), .B1(new_n588_), .B2(new_n572_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n794_), .A2(new_n799_), .A3(new_n596_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n548_), .B2(new_n543_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n800_), .B(KEYINPUT116), .C1(new_n548_), .C2(new_n543_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n662_), .B1(new_n786_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n504_), .A2(new_n807_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n786_), .B2(new_n805_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT118), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n780_), .A2(new_n781_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT117), .A3(new_n771_), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n780_), .A2(KEYINPUT117), .A3(new_n781_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n800_), .A2(new_n542_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n813_), .A2(new_n814_), .A3(KEYINPUT58), .A4(new_n815_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n670_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n809_), .C1(new_n786_), .C2(new_n805_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n808_), .A2(new_n811_), .A3(new_n820_), .A4(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n618_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n714_), .B1(new_n549_), .B2(new_n547_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n627_), .B2(new_n826_), .ZN(new_n827_));
  AND4_X1   g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n668_), .A4(new_n669_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n765_), .B1(new_n824_), .B2(new_n830_), .ZN(new_n831_));
  AOI211_X1 g630(.A(KEYINPUT119), .B(new_n829_), .C1(new_n823_), .C2(new_n618_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n764_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT120), .ZN(new_n834_));
  INV_X1    g633(.A(G113gat), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n836_), .B(new_n764_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n597_), .A4(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n824_), .A2(new_n830_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n764_), .B1(new_n840_), .B2(KEYINPUT59), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n764_), .A2(new_n840_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n839_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n833_), .B2(KEYINPUT59), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n844_), .A2(new_n597_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n838_), .B1(new_n845_), .B2(new_n835_), .ZN(G1340gat));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n844_), .B2(new_n551_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n849_));
  AOI21_X1  g648(.A(G120gat), .B1(new_n551_), .B2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n849_), .B2(G120gat), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n834_), .A2(new_n837_), .A3(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT122), .B1(new_n848_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n834_), .A2(new_n837_), .A3(new_n851_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n550_), .B(new_n843_), .C1(KEYINPUT59), .C2(new_n833_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n854_), .B(new_n855_), .C1(new_n856_), .C2(new_n847_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(G1341gat));
  AND3_X1   g657(.A1(new_n844_), .A2(G127gat), .A3(new_n628_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n834_), .A2(new_n628_), .A3(new_n837_), .ZN(new_n860_));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(KEYINPUT123), .A3(new_n861_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n859_), .B1(new_n864_), .B2(new_n865_), .ZN(G1342gat));
  INV_X1    g665(.A(G134gat), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n834_), .A2(new_n867_), .A3(new_n504_), .A4(new_n837_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n844_), .A2(new_n670_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1343gat));
  OR2_X1    g669(.A1(new_n831_), .A2(new_n832_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n647_), .A2(new_n394_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n686_), .A2(new_n634_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT124), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT124), .B(new_n873_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G141gat), .B1(new_n877_), .B2(new_n598_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n325_), .B(new_n597_), .C1(new_n874_), .C2(new_n876_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1344gat));
  OAI21_X1  g679(.A(G148gat), .B1(new_n877_), .B2(new_n550_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n326_), .B(new_n551_), .C1(new_n874_), .C2(new_n876_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1345gat));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n877_), .B2(new_n618_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n884_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n628_), .B(new_n886_), .C1(new_n874_), .C2(new_n876_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1346gat));
  OAI21_X1  g687(.A(G162gat), .B1(new_n877_), .B2(new_n627_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n662_), .A2(G162gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1347gat));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n739_), .A2(new_n647_), .A3(new_n638_), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n652_), .B(new_n894_), .C1(new_n824_), .C2(new_n830_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n895_), .A2(new_n597_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT22), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n893_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G169gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n210_), .B1(new_n896_), .B2(new_n893_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(new_n900_), .ZN(G1348gat));
  AOI21_X1  g700(.A(G176gat), .B1(new_n895_), .B2(new_n551_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n871_), .A2(new_n394_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n894_), .A2(new_n550_), .A3(new_n211_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(G1349gat));
  NOR2_X1   g704(.A1(new_n894_), .A2(new_n618_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n871_), .A2(new_n394_), .A3(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(G183gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n220_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n895_), .A2(new_n910_), .A3(new_n628_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n909_), .A2(KEYINPUT125), .A3(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1350gat));
  AOI21_X1  g715(.A(new_n218_), .B1(new_n895_), .B2(new_n670_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT126), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n895_), .A2(new_n221_), .A3(new_n504_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1351gat));
  AND3_X1   g719(.A1(new_n638_), .A2(new_n872_), .A3(new_n716_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n871_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n597_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n551_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G204gat), .ZN(G1353gat));
  OAI211_X1 g725(.A(new_n628_), .B(new_n921_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT63), .B(G211gat), .Z(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT127), .ZN(G1354gat));
  INV_X1    g730(.A(G218gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n922_), .A2(new_n932_), .A3(new_n504_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n922_), .A2(new_n670_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n933_), .B1(new_n935_), .B2(new_n932_), .ZN(G1355gat));
endmodule


