//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT77), .B(G43gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G99gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(G190gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n211_), .B(new_n212_), .C1(G183gat), .C2(G190gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(G169gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n217_), .A2(new_n218_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n211_), .A2(new_n212_), .ZN(new_n225_));
  INV_X1    g024(.A(G169gat), .ZN(new_n226_));
  INV_X1    g025(.A(G176gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(KEYINPUT24), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n230_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n216_), .B1(new_n224_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT30), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n207_), .B1(new_n234_), .B2(KEYINPUT78), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n232_), .B(KEYINPUT30), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n235_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n240_));
  INV_X1    g039(.A(G134gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G127gat), .ZN(new_n242_));
  INV_X1    g041(.A(G127gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G134gat), .ZN(new_n244_));
  INV_X1    g043(.A(G120gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G113gat), .ZN(new_n246_));
  INV_X1    g045(.A(G113gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G120gat), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n242_), .A2(new_n244_), .A3(new_n246_), .A4(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n242_), .A2(new_n244_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n240_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n242_), .A2(new_n244_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n246_), .A2(new_n248_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT80), .A3(new_n249_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT31), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(KEYINPUT31), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n259_), .A2(KEYINPUT79), .A3(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n239_), .B(new_n261_), .Z(new_n262_));
  XOR2_X1   g061(.A(G155gat), .B(G162gat), .Z(new_n263_));
  INV_X1    g062(.A(KEYINPUT81), .ZN(new_n264_));
  OAI22_X1  g063(.A1(new_n264_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT2), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n265_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(KEYINPUT3), .ZN(new_n271_));
  INV_X1    g070(.A(G141gat), .ZN(new_n272_));
  INV_X1    g071(.A(G148gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT3), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT81), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n271_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n263_), .B1(new_n270_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT82), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT82), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n280_), .B(new_n263_), .C1(new_n270_), .C2(new_n277_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n274_), .A2(new_n266_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n284_), .B1(KEYINPUT1), .B2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(KEYINPUT1), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n283_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n257_), .B1(new_n282_), .B2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n250_), .A2(new_n251_), .ZN(new_n291_));
  AOI211_X1 g090(.A(new_n288_), .B(new_n291_), .C1(new_n279_), .C2(new_n281_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT4), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G225gat), .A2(G233gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n281_), .ZN(new_n296_));
  AND3_X1   g095(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n275_), .A2(new_n272_), .A3(new_n273_), .A4(KEYINPUT81), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n271_), .A4(new_n265_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n280_), .B1(new_n301_), .B2(new_n263_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n289_), .B1(new_n296_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n258_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT4), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n293_), .A2(new_n295_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n291_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n282_), .A2(new_n289_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n295_), .B1(new_n304_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G1gat), .B(G29gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G57gat), .B(G85gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT98), .B1(new_n312_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n318_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT98), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n307_), .A2(new_n321_), .A3(new_n317_), .A4(new_n311_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n262_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(KEYINPUT84), .A2(G233gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(KEYINPUT84), .A2(G233gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(G228gat), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G211gat), .B(G218gat), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G197gat), .A2(G204gat), .ZN(new_n332_));
  OR2_X1    g131(.A1(KEYINPUT86), .A2(G197gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(KEYINPUT86), .A2(G197gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n335_), .B2(G204gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n331_), .B1(new_n336_), .B2(KEYINPUT21), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G204gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n333_), .A2(new_n339_), .A3(new_n334_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT21), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(G197gat), .B2(G204gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT87), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT87), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(new_n345_), .A3(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n330_), .A2(KEYINPUT21), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n336_), .B2(KEYINPUT88), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT88), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n339_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n350_), .B1(new_n351_), .B2(new_n332_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n338_), .A2(new_n347_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(KEYINPUT85), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n303_), .A2(KEYINPUT29), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n329_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n329_), .A3(new_n355_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT89), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n288_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G22gat), .B(G50gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n364_), .B(KEYINPUT28), .ZN(new_n369_));
  INV_X1    g168(.A(new_n367_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n361_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n357_), .A2(new_n358_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(new_n359_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n371_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT83), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n368_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n360_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n376_), .A2(new_n378_), .B1(new_n380_), .B2(new_n361_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n374_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT18), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT19), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n336_), .A2(KEYINPUT88), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n390_), .A2(KEYINPUT21), .A3(new_n330_), .A4(new_n352_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n344_), .A2(new_n346_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(new_n337_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n209_), .A2(KEYINPUT25), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n209_), .A2(KEYINPUT25), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n218_), .A2(KEYINPUT90), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n398_), .A3(new_n217_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n220_), .A2(new_n221_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n230_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT92), .B1(G183gat), .B2(G190gat), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n225_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT92), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n213_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n409_), .A3(new_n215_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n393_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n413_));
  INV_X1    g212(.A(new_n232_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(new_n353_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n389_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n413_), .B1(new_n393_), .B2(new_n232_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n399_), .A2(new_n401_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT91), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n230_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(new_n353_), .A3(new_n410_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n417_), .A2(new_n422_), .A3(new_n389_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n386_), .B1(new_n416_), .B2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n353_), .B1(new_n421_), .B2(new_n410_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT20), .B1(new_n393_), .B2(new_n232_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n388_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n417_), .A2(new_n422_), .A3(new_n389_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n386_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT27), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n425_), .A2(new_n426_), .A3(new_n388_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n389_), .B1(new_n417_), .B2(new_n422_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n386_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT27), .A3(new_n430_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n382_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n325_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n312_), .B2(new_n318_), .ZN(new_n443_));
  AOI211_X1 g242(.A(KEYINPUT33), .B(new_n317_), .C1(new_n307_), .C2(new_n311_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n304_), .A2(new_n309_), .A3(new_n295_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT4), .B1(new_n303_), .B2(new_n258_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n309_), .B1(new_n362_), .B2(new_n257_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n447_), .B1(new_n448_), .B2(KEYINPUT4), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n317_), .B(new_n446_), .C1(new_n449_), .C2(new_n295_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n424_), .A2(new_n430_), .A3(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT94), .B1(new_n445_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT32), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n386_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT97), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(KEYINPUT97), .B(new_n454_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n454_), .B(KEYINPUT95), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT96), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n460_), .A2(new_n427_), .A3(KEYINPUT96), .A4(new_n428_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n323_), .A2(new_n459_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n310_), .B1(new_n449_), .B2(new_n295_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT33), .B1(new_n467_), .B2(new_n317_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n312_), .A2(new_n442_), .A3(new_n318_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n424_), .A2(new_n430_), .A3(new_n450_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n452_), .A2(new_n466_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n382_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT99), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT99), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n477_), .A3(new_n382_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n382_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(new_n324_), .A3(new_n439_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n262_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n441_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G29gat), .B(G36gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT68), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G43gat), .B(G50gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G1gat), .B(G8gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT14), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT70), .B(G1gat), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n490_), .B1(new_n491_), .B2(G8gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT71), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G15gat), .B(G22gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(KEYINPUT72), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT72), .B1(new_n493_), .B2(new_n494_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n489_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n495_), .A3(new_n488_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n487_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n487_), .B(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n502_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n503_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n498_), .A2(new_n500_), .A3(new_n487_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n510_), .B2(new_n501_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G113gat), .B(G141gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT74), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G169gat), .B(G197gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n507_), .A2(new_n511_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(KEYINPUT75), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT75), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n483_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G85gat), .B(G92gat), .Z(new_n529_));
  NOR2_X1   g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n529_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT8), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(KEYINPUT9), .B2(new_n529_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(KEYINPUT10), .B(G99gat), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI221_X1 g340(.A(new_n538_), .B1(KEYINPUT9), .B2(new_n539_), .C1(G106gat), .C2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n537_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n487_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT35), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n487_), .B(KEYINPUT15), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n545_), .B(new_n550_), .C1(new_n551_), .C2(new_n543_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n548_), .A2(new_n549_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n537_), .A2(new_n542_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n505_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n553_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n545_), .A4(new_n550_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n554_), .A2(new_n563_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n557_), .B(KEYINPUT36), .Z(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT69), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n564_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n566_), .B1(new_n554_), .B2(new_n563_), .ZN(new_n572_));
  OAI211_X1 g371(.A(KEYINPUT69), .B(KEYINPUT37), .C1(new_n571_), .C2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n498_), .A2(new_n500_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(G231gat), .A3(G233gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n498_), .A2(new_n500_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G57gat), .B(G64gat), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n581_), .A2(KEYINPUT11), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(KEYINPUT11), .ZN(new_n583_));
  XOR2_X1   g382(.A(G71gat), .B(G78gat), .Z(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n583_), .A2(new_n584_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT73), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n580_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G127gat), .B(G155gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT16), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n577_), .A2(new_n588_), .A3(new_n579_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n590_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n594_), .A2(new_n595_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n590_), .B2(new_n597_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n575_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT13), .ZN(new_n604_));
  INV_X1    g403(.A(G230gat), .ZN(new_n605_));
  INV_X1    g404(.A(G233gat), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n537_), .A2(new_n542_), .A3(new_n587_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT64), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n543_), .A2(new_n587_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n608_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT12), .ZN(new_n615_));
  INV_X1    g414(.A(new_n587_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n560_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n615_), .B1(new_n560_), .B2(new_n616_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n614_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G120gat), .B(G148gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT65), .B(KEYINPUT5), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n612_), .A2(new_n620_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n612_), .B2(new_n620_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n604_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n629_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(KEYINPUT13), .A3(new_n627_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT66), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n603_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n528_), .A2(new_n635_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n636_), .A2(new_n324_), .A3(new_n491_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT38), .Z(new_n638_));
  INV_X1    g437(.A(new_n567_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n633_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n518_), .A2(new_n520_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n601_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n382_), .A2(new_n323_), .A3(new_n438_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n475_), .B2(KEYINPUT99), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n262_), .B1(new_n645_), .B2(new_n478_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n639_), .B(new_n643_), .C1(new_n646_), .C2(new_n441_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n324_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n638_), .A2(new_n648_), .ZN(G1324gat));
  OR3_X1    g448(.A1(new_n636_), .A2(G8gat), .A3(new_n439_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n651_), .B(G8gat), .C1(new_n647_), .C2(new_n439_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n483_), .A2(new_n567_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(new_n438_), .A3(new_n643_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n651_), .B1(new_n655_), .B2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n650_), .B1(new_n653_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT101), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n650_), .B(new_n659_), .C1(new_n653_), .C2(new_n656_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n658_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  OAI21_X1  g463(.A(G15gat), .B1(new_n647_), .B2(new_n482_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n482_), .A2(G15gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n636_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT103), .ZN(G1326gat));
  OAI21_X1  g469(.A(G22gat), .B1(new_n647_), .B2(new_n382_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT42), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n382_), .A2(G22gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n636_), .B2(new_n673_), .ZN(G1327gat));
  NAND2_X1  g473(.A1(new_n601_), .A2(new_n567_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n633_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n528_), .A2(new_n676_), .ZN(new_n677_));
  OR3_X1    g476(.A1(new_n677_), .A2(G29gat), .A3(new_n324_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n574_), .B(KEYINPUT104), .Z(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n483_), .B2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n575_), .A2(KEYINPUT43), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT105), .B1(new_n483_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n684_), .B(new_n681_), .C1(new_n646_), .C2(new_n441_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n680_), .A2(new_n683_), .A3(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n642_), .A2(new_n602_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n686_), .A2(new_n691_), .A3(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(KEYINPUT107), .A3(new_n323_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G29gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT107), .B1(new_n693_), .B2(new_n323_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n678_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n528_), .A2(new_n698_), .A3(new_n438_), .A4(new_n676_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT45), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n439_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n698_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n700_), .B(KEYINPUT46), .C1(new_n701_), .C2(new_n698_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  NAND2_X1  g505(.A1(new_n262_), .A2(G43gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT108), .B(G43gat), .Z(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n677_), .B2(new_n482_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n708_), .A2(KEYINPUT47), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT47), .B1(new_n708_), .B2(new_n711_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1330gat));
  INV_X1    g513(.A(new_n677_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G50gat), .B1(new_n715_), .B2(new_n479_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n479_), .A2(G50gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n693_), .B2(new_n717_), .ZN(G1331gat));
  AOI21_X1  g517(.A(new_n601_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n634_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n654_), .A2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n324_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n483_), .A2(new_n641_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n723_), .A2(new_n602_), .A3(new_n633_), .A4(new_n575_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n324_), .A2(G57gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n724_), .B2(new_n725_), .ZN(G1332gat));
  OAI21_X1  g525(.A(G64gat), .B1(new_n721_), .B2(new_n439_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT48), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n439_), .A2(G64gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n724_), .B2(new_n729_), .ZN(G1333gat));
  OAI21_X1  g529(.A(G71gat), .B1(new_n721_), .B2(new_n482_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT49), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n482_), .A2(G71gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n724_), .B2(new_n733_), .ZN(G1334gat));
  NAND3_X1  g533(.A1(new_n654_), .A2(new_n479_), .A3(new_n720_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(G78gat), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n735_), .B2(G78gat), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n382_), .A2(G78gat), .ZN(new_n740_));
  OAI22_X1  g539(.A1(new_n738_), .A2(new_n739_), .B1(new_n724_), .B2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT109), .Z(G1335gat));
  INV_X1    g541(.A(G85gat), .ZN(new_n743_));
  INV_X1    g542(.A(new_n634_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(new_n675_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n723_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n743_), .B1(new_n746_), .B2(new_n324_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT110), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n640_), .A2(new_n602_), .A3(new_n641_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n686_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n324_), .A2(new_n743_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(G1336gat));
  NOR3_X1   g551(.A1(new_n746_), .A2(G92gat), .A3(new_n439_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n686_), .A2(new_n438_), .A3(new_n749_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(G92gat), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT111), .Z(G1337gat));
  AND4_X1   g555(.A1(new_n262_), .A2(new_n723_), .A3(new_n540_), .A4(new_n745_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT112), .Z(new_n758_));
  NAND2_X1  g557(.A1(new_n750_), .A2(new_n262_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(G99gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(KEYINPUT113), .A3(KEYINPUT51), .ZN(new_n762_));
  NAND2_X1  g561(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n758_), .A2(new_n760_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1338gat));
  XNOR2_X1  g564(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n686_), .A2(new_n479_), .A3(new_n749_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G106gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT52), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  OR3_X1    g571(.A1(new_n746_), .A2(G106gat), .A3(new_n382_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n766_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n767_), .A2(new_n770_), .A3(G106gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n770_), .B1(new_n767_), .B2(G106gat), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n773_), .B(new_n766_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n774_), .A2(new_n778_), .ZN(G1339gat));
  INV_X1    g578(.A(KEYINPUT58), .ZN(new_n780_));
  INV_X1    g579(.A(new_n619_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n613_), .B1(new_n781_), .B2(new_n617_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT115), .B1(new_n782_), .B2(KEYINPUT55), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n620_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n618_), .A2(new_n619_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n607_), .B1(new_n787_), .B2(new_n610_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n782_), .A2(KEYINPUT55), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n783_), .A2(new_n786_), .A3(new_n788_), .A4(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n625_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n625_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n508_), .B1(new_n502_), .B2(new_n509_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT116), .B1(new_n795_), .B2(new_n516_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n503_), .B1(new_n510_), .B2(new_n501_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n515_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n502_), .A2(new_n508_), .A3(new_n506_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n796_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(new_n518_), .A3(new_n627_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n780_), .B1(new_n794_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n790_), .A2(new_n625_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n791_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n801_), .A2(new_n518_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(KEYINPUT58), .A4(new_n627_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n803_), .A2(new_n809_), .A3(new_n574_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n627_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n806_), .B2(new_n791_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n631_), .A2(new_n627_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n801_), .A2(new_n813_), .A3(new_n518_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n639_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT57), .B(new_n639_), .C1(new_n812_), .C2(new_n814_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n810_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n601_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT37), .B1(new_n567_), .B2(KEYINPUT69), .ZN(new_n822_));
  INV_X1    g621(.A(new_n573_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n633_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(new_n719_), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n824_), .B2(new_n719_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n821_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n440_), .A2(new_n482_), .A3(new_n324_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n818_), .B(KEYINPUT118), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n810_), .A2(new_n819_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n601_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n829_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n837_), .A2(new_n832_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n833_), .B1(new_n838_), .B2(new_n831_), .ZN(new_n839_));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839_), .B2(new_n527_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n247_), .A3(new_n641_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1340gat));
  OAI21_X1  g641(.A(G120gat), .B1(new_n839_), .B2(new_n744_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n245_), .B1(new_n640_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n838_), .B(new_n844_), .C1(KEYINPUT60), .C2(new_n245_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n839_), .B2(new_n601_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n838_), .A2(new_n243_), .A3(new_n602_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1342gat));
  OAI21_X1  g648(.A(G134gat), .B1(new_n839_), .B2(new_n575_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n838_), .A2(new_n241_), .A3(new_n567_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1343gat));
  NOR4_X1   g651(.A1(new_n262_), .A2(new_n382_), .A3(new_n324_), .A4(new_n438_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n837_), .A2(KEYINPUT119), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT119), .B1(new_n837_), .B2(new_n853_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n641_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g656(.A(new_n634_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g658(.A(new_n602_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1346gat));
  OR2_X1    g661(.A1(new_n854_), .A2(new_n855_), .ZN(new_n863_));
  INV_X1    g662(.A(G162gat), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n679_), .A2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n567_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n863_), .A2(new_n865_), .B1(new_n866_), .B2(new_n864_), .ZN(G1347gat));
  NOR2_X1   g666(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n226_), .B1(KEYINPUT122), .B2(KEYINPUT62), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n828_), .B1(new_n820_), .B2(new_n601_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n641_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n325_), .A2(new_n439_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT120), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n382_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n870_), .A2(new_n871_), .A3(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n869_), .B1(new_n876_), .B2(KEYINPUT121), .ZN(new_n877_));
  INV_X1    g676(.A(new_n875_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n830_), .A2(new_n641_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n868_), .B1(new_n877_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n876_), .A2(KEYINPUT121), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n880_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n868_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n869_), .A4(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT22), .B(G169gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n876_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n882_), .A2(new_n886_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT123), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n882_), .A2(new_n886_), .A3(new_n891_), .A4(new_n888_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1348gat));
  AOI21_X1  g692(.A(new_n479_), .B1(new_n836_), .B2(new_n829_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n873_), .A2(new_n744_), .A3(new_n227_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n830_), .A2(new_n633_), .A3(new_n878_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n894_), .A2(new_n895_), .B1(new_n896_), .B2(new_n227_), .ZN(G1349gat));
  NAND2_X1  g696(.A1(new_n830_), .A2(new_n878_), .ZN(new_n898_));
  AOI211_X1 g697(.A(new_n601_), .B(new_n898_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n894_), .A2(new_n602_), .A3(new_n874_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n900_), .A2(KEYINPUT124), .ZN(new_n901_));
  AOI21_X1  g700(.A(G183gat), .B1(new_n900_), .B2(KEYINPUT124), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n901_), .B2(new_n902_), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n898_), .B2(new_n575_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n567_), .A2(new_n217_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n898_), .B2(new_n905_), .ZN(G1351gat));
  NOR4_X1   g705(.A1(new_n262_), .A2(new_n382_), .A3(new_n439_), .A4(new_n323_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n837_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n641_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g709(.A1(new_n837_), .A2(new_n907_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n744_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n339_), .ZN(G1353gat));
  AOI21_X1  g712(.A(new_n601_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT125), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n908_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n916_), .B(new_n917_), .Z(G1354gat));
  NOR3_X1   g717(.A1(new_n911_), .A2(KEYINPUT126), .A3(new_n639_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(G218gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT126), .B1(new_n911_), .B2(new_n639_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n574_), .A2(G218gat), .ZN(new_n922_));
  XOR2_X1   g721(.A(new_n922_), .B(KEYINPUT127), .Z(new_n923_));
  AOI22_X1  g722(.A1(new_n920_), .A2(new_n921_), .B1(new_n908_), .B2(new_n923_), .ZN(G1355gat));
endmodule


