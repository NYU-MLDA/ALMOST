//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n959_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT10), .B(G99gat), .Z(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G85gat), .B(G92gat), .Z(new_n208_));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT64), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(KEYINPUT64), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n207_), .B(new_n212_), .C1(new_n213_), .C2(new_n210_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n204_), .A2(KEYINPUT65), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT7), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n215_), .B1(new_n222_), .B2(new_n208_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n208_), .A2(new_n215_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n224_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n214_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G71gat), .B(G78gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(KEYINPUT11), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT66), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n227_), .B(new_n232_), .C1(KEYINPUT11), .C2(new_n228_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n230_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n231_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT12), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT67), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n226_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n237_), .A2(KEYINPUT67), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G230gat), .A2(G233gat), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n226_), .A2(new_n236_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n226_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .A4(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n243_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n226_), .A2(new_n236_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n226_), .A2(new_n236_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G176gat), .B(G204gat), .Z(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT70), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G120gat), .B(G148gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT69), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n255_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n251_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(KEYINPUT13), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(KEYINPUT13), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n263_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G43gat), .B(G50gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(G29gat), .B(G36gat), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n268_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT78), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G15gat), .B(G22gat), .ZN(new_n273_));
  INV_X1    g072(.A(G1gat), .ZN(new_n274_));
  INV_X1    g073(.A(G8gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT14), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G1gat), .B(G8gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n272_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT15), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n271_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G229gat), .A2(G233gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT79), .ZN(new_n287_));
  INV_X1    g086(.A(new_n285_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n280_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n272_), .A2(new_n279_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT79), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n280_), .A2(new_n284_), .A3(new_n292_), .A4(new_n285_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n287_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G113gat), .B(G141gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G169gat), .B(G197gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n297_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n287_), .A2(new_n291_), .A3(new_n293_), .A4(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n266_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT21), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT96), .ZN(new_n309_));
  INV_X1    g108(.A(G197gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(new_n310_), .B2(G204gat), .ZN(new_n311_));
  INV_X1    g110(.A(G204gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(KEYINPUT96), .A3(G197gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(G204gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n308_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n311_), .A2(new_n313_), .A3(new_n307_), .A4(new_n314_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT97), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(G197gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n314_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT21), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n306_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n317_), .B1(new_n319_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT94), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G228gat), .A2(G233gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT95), .Z(new_n328_));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n330_));
  AND2_X1   g129(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT91), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n332_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n337_));
  OAI22_X1  g136(.A1(KEYINPUT91), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n338_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n330_), .B1(new_n337_), .B2(new_n343_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n333_), .A2(new_n336_), .B1(new_n340_), .B2(new_n339_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n331_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n345_), .A2(new_n348_), .A3(KEYINPUT92), .A4(new_n342_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n351_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT89), .B1(new_n352_), .B2(KEYINPUT1), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT90), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(KEYINPUT1), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT89), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT90), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(new_n356_), .A4(new_n351_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n352_), .A2(KEYINPUT1), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n359_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n333_), .A2(new_n339_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n329_), .B1(new_n355_), .B2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT96), .B1(new_n312_), .B2(G197gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n312_), .A2(G197gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n374_), .A2(KEYINPUT97), .A3(new_n307_), .A4(new_n313_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT97), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n318_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n323_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n316_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n326_), .B(new_n328_), .C1(new_n371_), .C2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n357_), .A2(new_n358_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n365_), .B1(new_n382_), .B2(new_n363_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n368_), .B1(new_n383_), .B2(new_n359_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n353_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT29), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n328_), .B1(new_n380_), .B2(KEYINPUT94), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n324_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n381_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n381_), .B2(new_n388_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n305_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n389_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n386_), .A2(new_n387_), .A3(new_n324_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n387_), .B1(new_n386_), .B2(new_n324_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n381_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n304_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n355_), .A2(new_n370_), .A3(new_n329_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G22gat), .B(G50gat), .Z(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n392_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n392_), .B2(new_n398_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT19), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT24), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G169gat), .A2(G176gat), .ZN(new_n409_));
  MUX2_X1   g208(.A(new_n408_), .B(KEYINPUT24), .S(new_n409_), .Z(new_n410_));
  INV_X1    g209(.A(KEYINPUT23), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(G183gat), .A3(G190gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G183gat), .A2(G190gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT82), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(G183gat), .A3(G190gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n412_), .B1(new_n417_), .B2(new_n411_), .ZN(new_n418_));
  INV_X1    g217(.A(G183gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n419_), .A2(KEYINPUT25), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT25), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(G183gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT26), .B(G190gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n410_), .A2(new_n418_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n407_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT22), .B(G169gat), .ZN(new_n429_));
  INV_X1    g228(.A(G176gat), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n417_), .A2(new_n433_), .A3(new_n411_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT23), .B1(new_n414_), .B2(new_n416_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT83), .B1(new_n413_), .B2(KEYINPUT23), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(G190gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n419_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n432_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n427_), .B1(new_n440_), .B2(KEYINPUT98), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT98), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n435_), .A2(new_n436_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n443_), .A2(new_n434_), .B1(new_n419_), .B2(new_n438_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n442_), .B1(new_n444_), .B2(new_n432_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n380_), .B1(new_n441_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n421_), .A2(G183gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT80), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n424_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n419_), .A2(KEYINPUT25), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n448_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT81), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT80), .B1(new_n420_), .B2(new_n422_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT81), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n424_), .A4(new_n449_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n437_), .A2(new_n410_), .A3(new_n453_), .A4(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n418_), .A2(new_n439_), .ZN(new_n458_));
  INV_X1    g257(.A(G169gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT22), .ZN(new_n460_));
  AOI21_X1  g259(.A(G176gat), .B1(new_n460_), .B2(KEYINPUT84), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(KEYINPUT84), .B2(new_n429_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n462_), .A3(new_n407_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n457_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT20), .B1(new_n464_), .B2(new_n324_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n406_), .B1(new_n446_), .B2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G8gat), .B(G36gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT18), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G64gat), .B(G92gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n441_), .A2(new_n445_), .A3(new_n380_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n406_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n473_), .B1(new_n464_), .B2(new_n324_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n466_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n470_), .B1(new_n466_), .B2(new_n475_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(KEYINPUT99), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT99), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n466_), .A2(new_n479_), .A3(new_n470_), .A4(new_n475_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT27), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n476_), .A2(KEYINPUT27), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n470_), .B(KEYINPUT101), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n437_), .A2(new_n439_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(KEYINPUT98), .A3(new_n431_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n426_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n440_), .A2(KEYINPUT98), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n324_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n465_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n472_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n380_), .B(new_n426_), .C1(new_n444_), .C2(new_n432_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n474_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n406_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n485_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n484_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G127gat), .B(G134gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G113gat), .B(G120gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n500_), .A2(new_n502_), .A3(KEYINPUT87), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n499_), .A2(new_n501_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT86), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n499_), .A2(new_n501_), .A3(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n503_), .A2(new_n507_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n355_), .A2(new_n370_), .A3(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(KEYINPUT4), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G225gat), .A2(G233gat), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n511_), .B1(new_n355_), .B2(new_n370_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G1gat), .B(G29gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT0), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(G57gat), .Z(new_n526_));
  INV_X1    g325(.A(G85gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n526_), .B(G85gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n521_), .A2(new_n522_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G71gat), .B(G99gat), .ZN(new_n533_));
  INV_X1    g332(.A(G43gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G227gat), .A2(G233gat), .ZN(new_n536_));
  INV_X1    g335(.A(G15gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n535_), .B(new_n538_), .Z(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT85), .B(KEYINPUT30), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n464_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n464_), .A2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n540_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(new_n542_), .A3(new_n539_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n545_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n511_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n545_), .A2(new_n547_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT31), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n545_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n512_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n532_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n404_), .A2(new_n483_), .A3(new_n498_), .A4(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT102), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n497_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n560_), .A2(new_n404_), .A3(KEYINPUT102), .A4(new_n556_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n392_), .A2(new_n398_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n401_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n392_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n532_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n521_), .A2(KEYINPUT33), .A3(new_n522_), .A4(new_n530_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n513_), .A2(G225gat), .A3(G233gat), .A4(new_n515_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n513_), .A2(KEYINPUT4), .A3(new_n515_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n517_), .B1(new_n513_), .B2(KEYINPUT4), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n528_), .B(new_n568_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n531_), .A2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n478_), .A2(new_n572_), .A3(new_n480_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n470_), .A2(KEYINPUT32), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n466_), .A2(new_n475_), .A3(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT100), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT100), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n466_), .A2(new_n581_), .A3(new_n475_), .A4(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n575_), .A2(new_n584_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n560_), .A2(new_n566_), .B1(new_n585_), .B2(new_n404_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n551_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n555_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n587_), .A2(new_n588_), .A3(KEYINPUT88), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT88), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n559_), .B(new_n561_), .C1(new_n586_), .C2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n303_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n223_), .A2(new_n225_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n271_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n214_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT34), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT35), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n226_), .A2(new_n282_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n605_), .A2(KEYINPUT72), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(KEYINPUT72), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n604_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n601_), .A2(new_n602_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G190gat), .B(G218gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT73), .ZN(new_n612_));
  XOR2_X1   g411(.A(G134gat), .B(G162gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n605_), .B(KEYINPUT72), .ZN(new_n617_));
  INV_X1    g416(.A(new_n609_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n604_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n610_), .A2(new_n616_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n614_), .B(new_n615_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n610_), .B2(new_n619_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n595_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n610_), .A2(new_n616_), .A3(new_n619_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n619_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n618_), .B1(new_n617_), .B2(new_n604_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT37), .B(new_n624_), .C1(new_n627_), .C2(new_n621_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n236_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n279_), .B(KEYINPUT74), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G183gat), .B(G211gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT76), .ZN(new_n635_));
  XOR2_X1   g434(.A(G127gat), .B(G155gat), .Z(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT77), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n637_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT17), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n633_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT17), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n633_), .B1(new_n643_), .B2(new_n640_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n629_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n594_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n274_), .A3(new_n532_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n620_), .A2(new_n622_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n593_), .A2(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n266_), .A2(new_n302_), .A3(new_n645_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n532_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n650_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1324gat));
  INV_X1    g460(.A(new_n560_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n655_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT105), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n655_), .A2(new_n665_), .A3(new_n662_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n664_), .A2(G8gat), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT39), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n664_), .A2(new_n669_), .A3(G8gat), .A4(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n647_), .A2(new_n275_), .A3(new_n662_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(KEYINPUT40), .A3(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  INV_X1    g476(.A(new_n592_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G15gat), .B1(new_n656_), .B2(new_n678_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n679_), .A2(KEYINPUT41), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(KEYINPUT41), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n647_), .A2(new_n537_), .A3(new_n592_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n680_), .A2(new_n681_), .A3(new_n682_), .ZN(G1326gat));
  INV_X1    g482(.A(G22gat), .ZN(new_n684_));
  INV_X1    g483(.A(new_n404_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n655_), .B2(new_n685_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT42), .Z(new_n687_));
  NAND3_X1  g486(.A1(new_n647_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(new_n645_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n652_), .A2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n594_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G29gat), .B1(new_n692_), .B2(new_n532_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n303_), .A2(new_n645_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n593_), .A2(new_n695_), .A3(new_n629_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n593_), .B2(new_n629_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(KEYINPUT106), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n593_), .A2(new_n699_), .A3(new_n695_), .A4(new_n629_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n694_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(KEYINPUT44), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n701_), .B2(KEYINPUT44), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n698_), .A2(new_n700_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n694_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n711_), .A2(G29gat), .A3(new_n532_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n693_), .B1(new_n706_), .B2(new_n712_), .ZN(G1328gat));
  XOR2_X1   g512(.A(KEYINPUT108), .B(KEYINPUT46), .Z(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n560_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n560_), .A2(G36gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n594_), .A2(new_n691_), .A3(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT45), .Z(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n715_), .B1(new_n718_), .B2(new_n722_), .ZN(new_n723_));
  AOI211_X1 g522(.A(new_n721_), .B(new_n714_), .C1(new_n717_), .C2(G36gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  AOI21_X1  g524(.A(G43gat), .B1(new_n692_), .B2(new_n592_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n587_), .A2(new_n588_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n711_), .A2(G43gat), .A3(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n727_), .B1(new_n705_), .B2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n732_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n727_), .B(new_n734_), .C1(new_n705_), .C2(new_n730_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1330gat));
  AOI21_X1  g535(.A(G50gat), .B1(new_n692_), .B2(new_n685_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n711_), .A2(G50gat), .A3(new_n685_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n706_), .B2(new_n738_), .ZN(G1331gat));
  AND3_X1   g538(.A1(new_n593_), .A2(new_n302_), .A3(new_n266_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n646_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G57gat), .B1(new_n741_), .B2(new_n532_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n645_), .A2(new_n301_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n653_), .A2(new_n266_), .A3(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n532_), .A2(new_n745_), .A3(G57gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n745_), .B2(G57gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n742_), .B1(new_n744_), .B2(new_n747_), .ZN(G1332gat));
  INV_X1    g547(.A(G64gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n744_), .B2(new_n662_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n741_), .A2(new_n749_), .A3(new_n662_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT111), .ZN(G1333gat));
  INV_X1    g554(.A(G71gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n744_), .B2(new_n592_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT49), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n741_), .A2(new_n756_), .A3(new_n592_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1334gat));
  INV_X1    g559(.A(G78gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n744_), .B2(new_n685_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n404_), .A2(G78gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT113), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n741_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n767_), .ZN(G1335gat));
  AND2_X1   g567(.A1(new_n740_), .A2(new_n691_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G85gat), .B1(new_n769_), .B2(new_n532_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n266_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n771_), .A2(new_n301_), .A3(new_n690_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n707_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n707_), .A2(KEYINPUT114), .A3(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n532_), .A2(G85gat), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT115), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n770_), .B1(new_n777_), .B2(new_n779_), .ZN(G1336gat));
  INV_X1    g579(.A(G92gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n769_), .A2(new_n781_), .A3(new_n662_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n560_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n781_), .ZN(G1337gat));
  AOI21_X1  g583(.A(new_n678_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n785_));
  INV_X1    g584(.A(G99gat), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n769_), .A2(new_n206_), .A3(new_n729_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT116), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT51), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n789_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n791_), .B(new_n792_), .C1(new_n786_), .C2(new_n785_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(G1338gat));
  NAND3_X1  g593(.A1(new_n769_), .A2(new_n205_), .A3(new_n685_), .ZN(new_n795_));
  OAI21_X1  g594(.A(G106gat), .B1(new_n773_), .B2(new_n404_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n796_), .A2(KEYINPUT52), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(KEYINPUT52), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n795_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n795_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n729_), .A2(new_n532_), .A3(new_n404_), .A4(new_n560_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n805_), .A2(KEYINPUT119), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(KEYINPUT119), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT120), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT59), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n629_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n743_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n266_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n266_), .A2(new_n816_), .A3(KEYINPUT54), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n246_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n249_), .B1(new_n248_), .B2(new_n240_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n825_), .A2(KEYINPUT55), .A3(new_n243_), .A4(new_n242_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n242_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n244_), .A2(new_n245_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n247_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n824_), .A2(new_n826_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n258_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n251_), .A2(new_n258_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n285_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n280_), .A2(new_n284_), .A3(new_n288_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n297_), .A3(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n300_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n833_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n832_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n831_), .B1(new_n830_), .B2(new_n258_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n822_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n830_), .A2(new_n258_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT56), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n843_), .A2(KEYINPUT58), .A3(new_n832_), .A4(new_n838_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n841_), .A2(new_n629_), .A3(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n259_), .A2(new_n300_), .A3(new_n836_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n842_), .A2(new_n847_), .A3(KEYINPUT56), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n302_), .A2(new_n833_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT56), .B1(new_n842_), .B2(new_n847_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n846_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n652_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n845_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n842_), .A2(new_n847_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n831_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n651_), .B1(new_n859_), .B2(new_n846_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n856_), .B1(new_n860_), .B2(KEYINPUT57), .ZN(new_n861_));
  AND4_X1   g660(.A1(new_n856_), .A2(new_n852_), .A3(KEYINPUT57), .A4(new_n652_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n855_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n645_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n821_), .B1(new_n864_), .B2(KEYINPUT121), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT118), .B1(new_n853_), .B2(new_n854_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n860_), .A2(new_n856_), .A3(KEYINPUT57), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n690_), .B1(new_n868_), .B2(new_n855_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n814_), .B1(new_n865_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n819_), .A2(new_n820_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n864_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n875_), .B2(new_n809_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n804_), .B1(new_n872_), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n874_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n864_), .A2(KEYINPUT121), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n813_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n869_), .A2(new_n821_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT59), .B1(new_n881_), .B2(new_n808_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(KEYINPUT122), .A3(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n877_), .A2(new_n883_), .A3(new_n301_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G113gat), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n881_), .A2(new_n808_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  OR3_X1    g686(.A1(new_n887_), .A2(G113gat), .A3(new_n302_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n888_), .ZN(G1340gat));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n890_));
  INV_X1    g689(.A(G120gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n266_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n886_), .A2(new_n893_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n872_), .A2(new_n876_), .A3(new_n771_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n891_), .ZN(G1341gat));
  NAND3_X1  g695(.A1(new_n877_), .A2(new_n883_), .A3(new_n690_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G127gat), .ZN(new_n898_));
  OR3_X1    g697(.A1(new_n887_), .A2(G127gat), .A3(new_n645_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1342gat));
  NAND3_X1  g699(.A1(new_n877_), .A2(new_n883_), .A3(new_n629_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G134gat), .ZN(new_n902_));
  OR3_X1    g701(.A1(new_n887_), .A2(G134gat), .A3(new_n652_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1343gat));
  NOR2_X1   g703(.A1(new_n592_), .A2(new_n404_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n662_), .A2(new_n657_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n905_), .B(new_n906_), .C1(new_n869_), .C2(new_n821_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n302_), .ZN(new_n908_));
  XOR2_X1   g707(.A(new_n908_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n771_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(G148gat), .Z(G1345gat));
  XOR2_X1   g710(.A(KEYINPUT61), .B(G155gat), .Z(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT123), .B1(new_n907_), .B2(new_n645_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n905_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n874_), .B2(new_n864_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n915_), .A2(new_n916_), .A3(new_n690_), .A4(new_n906_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n913_), .A2(new_n917_), .A3(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n913_), .B2(new_n917_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n912_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n913_), .A2(new_n917_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT124), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n913_), .A2(new_n917_), .A3(new_n918_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n912_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n921_), .A2(new_n926_), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n907_), .B2(new_n815_), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n652_), .A2(G162gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n907_), .B2(new_n929_), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n560_), .A2(new_n532_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n592_), .A2(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT125), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n685_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n934_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT126), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n937_), .B(new_n934_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n939_), .A2(new_n429_), .A3(new_n301_), .ZN(new_n940_));
  OAI21_X1  g739(.A(G169gat), .B1(new_n935_), .B2(new_n302_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n941_), .A2(KEYINPUT62), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(KEYINPUT62), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n940_), .B1(new_n942_), .B2(new_n943_), .ZN(G1348gat));
  NAND2_X1  g743(.A1(new_n939_), .A2(new_n266_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n881_), .A2(new_n685_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n933_), .A2(new_n430_), .A3(new_n771_), .ZN(new_n947_));
  AOI22_X1  g746(.A1(new_n945_), .A2(new_n430_), .B1(new_n946_), .B2(new_n947_), .ZN(G1349gat));
  NOR2_X1   g747(.A1(new_n933_), .A2(new_n645_), .ZN(new_n949_));
  AOI21_X1  g748(.A(G183gat), .B1(new_n946_), .B2(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n645_), .A2(new_n423_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n939_), .B2(new_n951_), .ZN(G1350gat));
  NAND3_X1  g751(.A1(new_n939_), .A2(new_n651_), .A3(new_n424_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n815_), .B1(new_n936_), .B2(new_n938_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n438_), .B2(new_n954_), .ZN(G1351gat));
  NAND2_X1  g754(.A1(new_n915_), .A2(new_n931_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n956_), .A2(new_n302_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(new_n310_), .ZN(G1352gat));
  NOR2_X1   g757(.A1(new_n956_), .A2(new_n771_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(new_n312_), .ZN(G1353gat));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961_));
  INV_X1    g760(.A(new_n956_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n645_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n961_), .B1(new_n964_), .B2(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n965_), .ZN(new_n967_));
  NAND4_X1  g766(.A1(new_n962_), .A2(KEYINPUT127), .A3(new_n967_), .A4(new_n963_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n964_), .A2(new_n965_), .ZN(new_n969_));
  AND3_X1   g768(.A1(new_n966_), .A2(new_n968_), .A3(new_n969_), .ZN(G1354gat));
  OAI21_X1  g769(.A(G218gat), .B1(new_n956_), .B2(new_n815_), .ZN(new_n971_));
  OR2_X1    g770(.A1(new_n652_), .A2(G218gat), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n956_), .B2(new_n972_), .ZN(G1355gat));
endmodule


