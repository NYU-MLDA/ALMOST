//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT15), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n208_));
  OAI22_X1  g007(.A1(new_n208_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n209_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT68), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n218_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n213_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G92gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT8), .B1(new_n221_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  INV_X1    g027(.A(new_n226_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n215_), .A2(new_n217_), .A3(KEYINPUT65), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT65), .B1(new_n215_), .B2(new_n217_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n228_), .B(new_n229_), .C1(new_n232_), .C2(new_n213_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235_));
  OR2_X1    g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n224_), .A2(KEYINPUT9), .A3(new_n225_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n225_), .A2(KEYINPUT9), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n235_), .B1(new_n232_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n215_), .A2(new_n217_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n215_), .A2(new_n217_), .A3(KEYINPUT65), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(KEYINPUT66), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n243_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n207_), .B1(new_n234_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G232gat), .A2(G233gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n254_), .B(KEYINPUT34), .Z(new_n255_));
  INV_X1    g054(.A(KEYINPUT35), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT73), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n227_), .A2(new_n233_), .B1(new_n243_), .B2(new_n250_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(new_n205_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n253_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n244_), .A2(KEYINPUT68), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n208_), .A2(KEYINPUT7), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n208_), .A2(KEYINPUT7), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n211_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n264_), .A2(new_n267_), .A3(new_n268_), .A4(new_n209_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n228_), .B1(new_n269_), .B2(new_n229_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n229_), .A2(new_n228_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n213_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n248_), .B2(new_n272_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n232_), .A2(new_n235_), .A3(new_n242_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT66), .B1(new_n248_), .B2(new_n249_), .ZN(new_n275_));
  OAI22_X1  g074(.A1(new_n270_), .A2(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n205_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n258_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT72), .B1(new_n278_), .B2(new_n252_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n263_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n255_), .A2(new_n256_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n263_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G190gat), .B(G218gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G134gat), .B(G162gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n283_), .A2(KEYINPUT36), .A3(new_n284_), .A4(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(KEYINPUT36), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n283_), .A2(new_n284_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n289_), .ZN(new_n293_));
  AOI211_X1 g092(.A(KEYINPUT74), .B(new_n293_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n288_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT23), .ZN(new_n297_));
  INV_X1    g096(.A(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(KEYINPUT24), .A3(new_n301_), .ZN(new_n302_));
  OR3_X1    g101(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT81), .B(G183gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT25), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT82), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G190gat), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(KEYINPUT83), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(KEYINPUT83), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n308_), .A2(G190gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT25), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(G183gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .A4(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n297_), .B(new_n304_), .C1(new_n307_), .C2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n301_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(G169gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n320_), .A2(G176gat), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n318_), .B(G169gat), .C1(new_n319_), .C2(KEYINPUT22), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n317_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n296_), .B2(KEYINPUT23), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n297_), .B2(new_n324_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n305_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(G190gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n323_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n316_), .A2(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(KEYINPUT87), .B(G15gat), .Z(new_n331_));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n330_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G113gat), .B(G120gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n334_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G71gat), .B(G99gat), .ZN(new_n339_));
  INV_X1    g138(.A(G43gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT30), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT31), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n338_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n348_));
  INV_X1    g147(.A(G141gat), .ZN(new_n349_));
  INV_X1    g148(.A(G148gat), .ZN(new_n350_));
  OAI211_X1 g149(.A(KEYINPUT89), .B(new_n348_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  OR3_X1    g150(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT89), .B1(new_n349_), .B2(new_n350_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT2), .ZN(new_n356_));
  AOI211_X1 g155(.A(new_n346_), .B(new_n347_), .C1(new_n354_), .C2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G141gat), .B(G148gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n345_), .B1(new_n347_), .B2(KEYINPUT1), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n359_), .A2(KEYINPUT88), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n345_), .A2(KEYINPUT1), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n359_), .B2(KEYINPUT88), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n358_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT28), .ZN(new_n367_));
  XOR2_X1   g166(.A(G22gat), .B(G50gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT92), .Z(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n372_), .A2(KEYINPUT93), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT90), .B(G204gat), .ZN(new_n376_));
  INV_X1    g175(.A(G197gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT91), .Z(new_n379_));
  XOR2_X1   g178(.A(G211gat), .B(G218gat), .Z(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(KEYINPUT21), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n377_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT21), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(G197gat), .B2(G204gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n378_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n385_), .B1(new_n386_), .B2(KEYINPUT21), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n364_), .A2(new_n365_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G228gat), .A2(G233gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n369_), .A2(new_n372_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n374_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n393_), .B1(new_n374_), .B2(new_n394_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n388_), .A2(new_n330_), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n400_), .B(KEYINPUT95), .Z(new_n401_));
  INV_X1    g200(.A(KEYINPUT20), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT19), .ZN(new_n404_));
  XOR2_X1   g203(.A(KEYINPUT25), .B(G183gat), .Z(new_n405_));
  NAND2_X1  g204(.A1(new_n312_), .A2(new_n309_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n304_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(new_n326_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT94), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n297_), .B1(G183gat), .B2(G190gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT22), .B(G169gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n317_), .B1(new_n412_), .B2(new_n299_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  AOI211_X1 g214(.A(new_n402_), .B(new_n404_), .C1(new_n415_), .C2(new_n389_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n401_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n388_), .A2(new_n330_), .ZN(new_n418_));
  OAI211_X1 g217(.A(KEYINPUT20), .B(new_n418_), .C1(new_n415_), .C2(new_n389_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n404_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT18), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n417_), .A2(new_n420_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n425_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G85gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT0), .B(G57gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n431_), .B(new_n432_), .Z(new_n433_));
  NOR3_X1   g232(.A1(new_n357_), .A2(KEYINPUT96), .A3(new_n363_), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n434_), .B(new_n337_), .Z(new_n435_));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT97), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT98), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n433_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n337_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT99), .Z(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n437_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n435_), .A2(KEYINPUT4), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n440_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n426_), .A2(new_n429_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n435_), .A2(new_n437_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n439_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n433_), .B(new_n447_), .C1(new_n448_), .C2(new_n444_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT100), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n450_), .A2(KEYINPUT33), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(KEYINPUT33), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n446_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n425_), .A2(KEYINPUT32), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n421_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n404_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n408_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n402_), .B1(new_n389_), .B2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n456_), .B1(new_n401_), .B2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n419_), .A2(new_n404_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n455_), .B1(new_n461_), .B2(new_n454_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n447_), .B1(new_n448_), .B2(new_n444_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n433_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n465_), .A2(new_n449_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n462_), .A2(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n344_), .B(new_n399_), .C1(new_n453_), .C2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n426_), .A2(new_n429_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(new_n421_), .B2(new_n425_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n428_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n469_), .A2(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n344_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n374_), .A2(new_n394_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n393_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(new_n344_), .A3(new_n395_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n466_), .B(new_n473_), .C1(new_n476_), .C2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n295_), .B1(new_n468_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G230gat), .A2(G233gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n484_), .B(KEYINPUT64), .Z(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n488_));
  XOR2_X1   g287(.A(G71gat), .B(G78gat), .Z(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n488_), .A2(new_n489_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n260_), .A2(new_n492_), .B1(KEYINPUT69), .B2(KEYINPUT12), .ZN(new_n493_));
  INV_X1    g292(.A(new_n492_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n276_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n495_), .B1(new_n276_), .B2(new_n494_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n485_), .B(new_n493_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n485_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n260_), .A2(new_n492_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n276_), .A2(new_n494_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n499_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G120gat), .B(G148gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G176gat), .B(G204gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n498_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n507_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n511_), .B1(new_n514_), .B2(new_n512_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n207_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518_));
  INV_X1    g317(.A(G8gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G1gat), .B(G8gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT78), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n524_), .B(new_n526_), .C1(new_n523_), .C2(new_n277_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n523_), .B(new_n205_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT77), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n529_), .B2(new_n525_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT79), .B(KEYINPUT80), .Z(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n530_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n516_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G231gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n523_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(new_n492_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT75), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(KEYINPUT75), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G127gat), .B(G155gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT16), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G183gat), .B(G211gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT17), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT76), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n542_), .A2(new_n543_), .A3(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n547_), .A2(KEYINPUT17), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n541_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n538_), .A2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n483_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n466_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n202_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT101), .Z(new_n558_));
  AOI21_X1  g357(.A(new_n536_), .B1(new_n468_), .B2(new_n482_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n295_), .A2(KEYINPUT37), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n561_), .B(new_n288_), .C1(new_n292_), .C2(new_n294_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(new_n553_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n516_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n559_), .A2(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n567_), .A2(G1gat), .A3(new_n466_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT38), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(KEYINPUT38), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n558_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT102), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT102), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n558_), .A2(new_n573_), .A3(new_n569_), .A4(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(G1324gat));
  INV_X1    g374(.A(new_n567_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n473_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n519_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n555_), .A2(new_n577_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(G8gat), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n580_), .A2(KEYINPUT39), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(KEYINPUT39), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n578_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT40), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(G1325gat));
  INV_X1    g384(.A(G15gat), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n555_), .B2(new_n474_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT41), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n576_), .A2(new_n586_), .A3(new_n474_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(G1326gat));
  INV_X1    g389(.A(G22gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n398_), .B(KEYINPUT103), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n555_), .B2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n576_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(G1327gat));
  INV_X1    g396(.A(new_n295_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n553_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n559_), .A2(new_n516_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(G29gat), .B1(new_n601_), .B2(new_n556_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n468_), .A2(new_n482_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n563_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT43), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT43), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(new_n606_), .A3(new_n563_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n538_), .A2(new_n599_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT44), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT44), .ZN(new_n611_));
  INV_X1    g410(.A(new_n609_), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n611_), .B(new_n612_), .C1(new_n605_), .C2(new_n607_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n556_), .A2(G29gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n602_), .B1(new_n614_), .B2(new_n615_), .ZN(G1328gat));
  INV_X1    g415(.A(KEYINPUT105), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(KEYINPUT46), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n473_), .A2(G36gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n601_), .A2(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT45), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(KEYINPUT45), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n618_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n610_), .A2(new_n613_), .A3(new_n473_), .ZN(new_n624_));
  INV_X1    g423(.A(G36gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n623_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n617_), .A2(KEYINPUT46), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT106), .Z(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n623_), .B(new_n628_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1329gat));
  AOI21_X1  g431(.A(G43gat), .B1(new_n601_), .B2(new_n474_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n344_), .A2(new_n340_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n614_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT47), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(G1330gat));
  AOI21_X1  g436(.A(G50gat), .B1(new_n601_), .B2(new_n592_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n398_), .A2(G50gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n614_), .B2(new_n639_), .ZN(G1331gat));
  NOR3_X1   g439(.A1(new_n516_), .A2(new_n537_), .A3(new_n553_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n483_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n556_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G57gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n537_), .B1(new_n468_), .B2(new_n482_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n516_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n564_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n466_), .A2(G57gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n644_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT107), .Z(G1332gat));
  INV_X1    g450(.A(G64gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n642_), .B2(new_n577_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT48), .Z(new_n654_));
  INV_X1    g453(.A(new_n648_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n652_), .A3(new_n577_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1333gat));
  NAND2_X1  g456(.A1(new_n642_), .A2(new_n474_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(G71gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n344_), .A2(G71gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT109), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n648_), .B2(new_n663_), .ZN(G1334gat));
  INV_X1    g463(.A(G78gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n655_), .A2(new_n665_), .A3(new_n592_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n642_), .A2(new_n592_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G78gat), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(KEYINPUT50), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(KEYINPUT50), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT110), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(G1335gat));
  NOR2_X1   g472(.A1(new_n537_), .A2(new_n599_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n646_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT111), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n608_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n605_), .A2(KEYINPUT111), .A3(new_n607_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G85gat), .B1(new_n680_), .B2(new_n466_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n645_), .A2(new_n646_), .A3(new_n600_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n222_), .A3(new_n556_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1336gat));
  OAI21_X1  g484(.A(G92gat), .B1(new_n680_), .B2(new_n473_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n683_), .A2(new_n223_), .A3(new_n577_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1337gat));
  INV_X1    g487(.A(G99gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n679_), .B2(new_n474_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT51), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(KEYINPUT112), .ZN(new_n692_));
  AND4_X1   g491(.A1(new_n474_), .A2(new_n683_), .A3(new_n236_), .A4(new_n238_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n690_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1338gat));
  NOR2_X1   g495(.A1(new_n675_), .A2(new_n399_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT113), .ZN(new_n700_));
  OR3_X1    g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n237_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(new_n237_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(KEYINPUT52), .A3(new_n702_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n702_), .A2(KEYINPUT52), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n683_), .A2(new_n237_), .A3(new_n398_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT53), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT53), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n703_), .A2(new_n704_), .A3(new_n708_), .A4(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1339gat));
  NOR2_X1   g509(.A1(new_n577_), .A2(new_n466_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n476_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(KEYINPUT59), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT54), .B1(new_n565_), .B2(new_n537_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT54), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n564_), .A2(new_n715_), .A3(new_n536_), .A4(new_n516_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n527_), .B(new_n535_), .C1(new_n529_), .C2(new_n525_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n523_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n526_), .B1(new_n719_), .B2(new_n205_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n535_), .B1(new_n524_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n526_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n529_), .B2(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n718_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n511_), .A2(KEYINPUT115), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT115), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT56), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n493_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n499_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n495_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n733_), .B1(new_n260_), .B2(new_n492_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n276_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n736_), .A2(KEYINPUT55), .A3(new_n485_), .A4(new_n493_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n732_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n498_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT114), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n740_), .A2(new_n732_), .A3(new_n737_), .A4(KEYINPUT114), .ZN(new_n742_));
  INV_X1    g541(.A(new_n507_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n730_), .B1(new_n741_), .B2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n732_), .A3(new_n737_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n748_), .A2(KEYINPUT56), .A3(new_n743_), .A4(new_n742_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n745_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n536_), .A2(new_n509_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n729_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT116), .B1(new_n752_), .B2(new_n295_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n724_), .A2(new_n508_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n745_), .B2(new_n749_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n755_), .A2(KEYINPUT58), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n755_), .A2(KEYINPUT58), .B1(new_n560_), .B2(new_n562_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n753_), .A2(KEYINPUT57), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT116), .B(new_n759_), .C1(new_n752_), .C2(new_n295_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n599_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT118), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n717_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT118), .B(new_n599_), .C1(new_n758_), .C2(new_n760_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n713_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n753_), .A2(KEYINPUT57), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n757_), .A2(new_n756_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n760_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n758_), .A2(KEYINPUT117), .A3(new_n760_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n553_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n712_), .B1(new_n772_), .B2(new_n717_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT59), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n765_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G113gat), .B1(new_n775_), .B2(new_n536_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n773_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n536_), .A2(G113gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(G1340gat));
  INV_X1    g578(.A(G120gat), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n765_), .B(new_n646_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(KEYINPUT119), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(KEYINPUT119), .B2(new_n781_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n516_), .B2(KEYINPUT60), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n773_), .B(new_n784_), .C1(KEYINPUT60), .C2(new_n780_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1341gat));
  OAI21_X1  g585(.A(G127gat), .B1(new_n775_), .B2(new_n553_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n553_), .A2(G127gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n777_), .B2(new_n788_), .ZN(G1342gat));
  OAI211_X1 g588(.A(new_n765_), .B(new_n563_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G134gat), .ZN(new_n791_));
  INV_X1    g590(.A(G134gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n773_), .A2(new_n792_), .A3(new_n295_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n791_), .A2(KEYINPUT120), .A3(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1343gat));
  XNOR2_X1  g597(.A(KEYINPUT122), .B(G141gat), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n772_), .A2(new_n717_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n481_), .A3(new_n711_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT121), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n480_), .B1(new_n772_), .B2(new_n717_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n711_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n799_), .B1(new_n806_), .B2(new_n537_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n799_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n536_), .B(new_n808_), .C1(new_n802_), .C2(new_n805_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n807_), .A2(new_n809_), .ZN(G1344gat));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n646_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G148gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n350_), .A3(new_n646_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1345gat));
  NAND2_X1  g613(.A1(new_n806_), .A2(new_n599_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT61), .B(G155gat), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n816_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n806_), .A2(new_n599_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1346gat));
  INV_X1    g619(.A(G162gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n806_), .A2(new_n821_), .A3(new_n295_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n563_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n802_), .B2(new_n805_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n821_), .B2(new_n824_), .ZN(G1347gat));
  NOR2_X1   g624(.A1(new_n473_), .A2(new_n556_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n474_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(new_n592_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n537_), .B(new_n828_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G169gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n768_), .A2(new_n553_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT118), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n761_), .A2(new_n762_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n717_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(new_n412_), .A3(new_n537_), .A4(new_n828_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n830_), .A2(KEYINPUT62), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n829_), .A2(new_n837_), .A3(G169gat), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT123), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n836_), .A2(new_n841_), .A3(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1348gat));
  AND2_X1   g642(.A1(new_n834_), .A2(new_n828_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G176gat), .B1(new_n844_), .B2(new_n646_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n599_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n846_), .A2(new_n771_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n398_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n827_), .A2(new_n299_), .A3(new_n516_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n845_), .B1(new_n848_), .B2(new_n849_), .ZN(G1349gat));
  NOR2_X1   g649(.A1(new_n827_), .A2(new_n553_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n848_), .A2(KEYINPUT124), .A3(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n599_), .A2(new_n405_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n856_), .A2(new_n305_), .B1(new_n844_), .B2(new_n858_), .ZN(G1350gat));
  NAND2_X1  g658(.A1(new_n844_), .A2(new_n563_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G190gat), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n598_), .A2(new_n406_), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT125), .Z(new_n863_));
  NAND2_X1  g662(.A1(new_n844_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n861_), .A2(new_n864_), .ZN(G1351gat));
  NAND3_X1  g664(.A1(new_n800_), .A2(new_n481_), .A3(new_n826_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT126), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n803_), .A2(KEYINPUT126), .A3(new_n826_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G197gat), .B1(new_n870_), .B2(new_n537_), .ZN(new_n871_));
  AOI211_X1 g670(.A(new_n377_), .B(new_n536_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1352gat));
  INV_X1    g672(.A(new_n376_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n803_), .A2(KEYINPUT126), .A3(new_n826_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT126), .B1(new_n803_), .B2(new_n826_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n874_), .B(new_n646_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n516_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(G204gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(G1353gat));
  XOR2_X1   g679(.A(KEYINPUT63), .B(G211gat), .Z(new_n881_));
  OAI211_X1 g680(.A(new_n599_), .B(new_n881_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n553_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n883_));
  OR2_X1    g682(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(G1354gat));
  INV_X1    g685(.A(G218gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n870_), .A2(new_n887_), .A3(new_n295_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n823_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n887_), .B2(new_n889_), .ZN(G1355gat));
endmodule


