//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(KEYINPUT36), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G232gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT34), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT10), .B(G99gat), .Z(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G85gat), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  OR3_X1    g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT9), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n213_), .A2(new_n216_), .A3(new_n219_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n229_), .A2(new_n222_), .A3(new_n223_), .A4(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n212_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n231_), .B2(new_n212_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n225_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G43gat), .B(G50gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(G29gat), .B(G36gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT69), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n238_), .B(KEYINPUT15), .Z(new_n241_));
  NOR3_X1   g040(.A1(new_n233_), .A2(new_n234_), .A3(KEYINPUT66), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n231_), .A2(new_n212_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT8), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n231_), .A2(new_n232_), .A3(new_n212_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n243_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n225_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n211_), .A2(KEYINPUT35), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(KEYINPUT35), .B(new_n211_), .C1(new_n240_), .C2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n239_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n211_), .A2(KEYINPUT35), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(new_n250_), .A4(new_n249_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n209_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n252_), .A2(new_n256_), .A3(KEYINPUT72), .A4(new_n208_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n206_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(KEYINPUT36), .A3(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n259_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT37), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G15gat), .B(G22gat), .ZN(new_n265_));
  INV_X1    g064(.A(G1gat), .ZN(new_n266_));
  INV_X1    g065(.A(G8gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT14), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G1gat), .B(G8gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G231gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G57gat), .ZN(new_n274_));
  INV_X1    g073(.A(G64gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G57gat), .A2(G64gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT11), .ZN(new_n279_));
  XOR2_X1   g078(.A(G71gat), .B(G78gat), .Z(new_n280_));
  OR2_X1    g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT11), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n276_), .A2(new_n282_), .A3(new_n277_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n273_), .B(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G183gat), .B(G211gat), .Z(new_n288_));
  XNOR2_X1  g087(.A(G127gat), .B(G155gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT17), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n287_), .A2(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n292_), .A2(KEYINPUT17), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n287_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n264_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n285_), .A2(KEYINPUT12), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n248_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n235_), .A2(new_n285_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT12), .B1(new_n235_), .B2(new_n285_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n301_), .A2(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G230gat), .A2(G233gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n248_), .A2(KEYINPUT67), .A3(new_n300_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .A4(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n225_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT66), .B1(new_n233_), .B2(new_n234_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n245_), .A2(new_n243_), .A3(new_n246_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n285_), .A2(KEYINPUT12), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n302_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n304_), .A2(new_n303_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n308_), .A2(new_n315_), .A3(new_n307_), .A4(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT68), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n309_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n235_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT65), .B1(new_n320_), .B2(new_n286_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n307_), .B1(new_n321_), .B2(new_n303_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(new_n303_), .B2(new_n321_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G120gat), .B(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(G204gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT5), .B(G176gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n319_), .A2(new_n323_), .A3(new_n329_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n331_), .A2(KEYINPUT13), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT13), .B1(new_n331_), .B2(new_n332_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT22), .B(G169gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n338_), .A2(KEYINPUT78), .ZN(new_n339_));
  INV_X1    g138(.A(G169gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT78), .B1(new_n340_), .B2(KEYINPUT22), .ZN(new_n341_));
  INV_X1    g140(.A(G176gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n337_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(G183gat), .B2(G190gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT79), .ZN(new_n347_));
  INV_X1    g146(.A(G183gat), .ZN(new_n348_));
  INV_X1    g147(.A(G190gat), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n348_), .A2(new_n349_), .A3(KEYINPUT23), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT77), .B(G190gat), .Z(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n348_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT80), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n352_), .A2(new_n357_), .A3(new_n354_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n344_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n348_), .A2(KEYINPUT25), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n360_), .A2(KEYINPUT76), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(KEYINPUT76), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n361_), .A2(new_n362_), .B1(new_n363_), .B2(G183gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT26), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n349_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n353_), .B2(new_n365_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n350_), .A2(new_n346_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n340_), .A2(new_n342_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n371_), .A2(KEYINPUT24), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(KEYINPUT24), .A3(new_n337_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n368_), .A2(new_n370_), .A3(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n359_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G71gat), .B(G99gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G43gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n376_), .B(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G113gat), .B(G120gat), .Z(new_n380_));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n381_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT30), .B(G15gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT81), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT31), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n386_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n379_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(new_n218_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT18), .B(G64gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT32), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G197gat), .B(G204gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT85), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n326_), .A2(G197gat), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n399_), .B(KEYINPUT21), .C1(KEYINPUT85), .C2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT86), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G211gat), .B(G218gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT21), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n405_), .B2(new_n398_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n398_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n359_), .B2(new_n375_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT20), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n370_), .B1(G183gat), .B2(G190gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n338_), .A2(new_n342_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n337_), .A3(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT26), .B(G190gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n363_), .A2(G183gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n360_), .A3(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n352_), .A2(new_n374_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n412_), .B1(new_n413_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n411_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT19), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(KEYINPUT92), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT20), .B1(new_n413_), .B2(new_n422_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n359_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n375_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n413_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n426_), .B(KEYINPUT89), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n426_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n411_), .B2(new_n423_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(KEYINPUT92), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n397_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G155gat), .B(G162gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT83), .ZN(new_n443_));
  OR2_X1    g242(.A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(new_n444_));
  NAND2_X1  g243(.A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n444_), .A2(new_n445_), .B1(G141gat), .B2(G148gat), .ZN(new_n446_));
  INV_X1    g245(.A(G141gat), .ZN(new_n447_));
  INV_X1    g246(.A(G148gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(KEYINPUT3), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G141gat), .A2(G148gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n446_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n443_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(G155gat), .A2(G162gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n457_), .B1(KEYINPUT1), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n459_), .B1(KEYINPUT1), .B2(new_n458_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n453_), .A3(new_n449_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n456_), .A2(new_n461_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT90), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n456_), .A2(new_n461_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(new_n384_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT4), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n463_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n462_), .A2(KEYINPUT90), .A3(KEYINPUT4), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G225gat), .A2(G233gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n465_), .A2(new_n462_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n471_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G1gat), .B(G29gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(new_n217_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT0), .B(G57gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n472_), .A2(new_n475_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n470_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n482_), .B2(new_n474_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n433_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n410_), .A2(new_n359_), .A3(new_n375_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n428_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n411_), .A2(new_n437_), .A3(new_n423_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n397_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n482_), .A2(new_n474_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n492_), .B2(new_n480_), .ZN(new_n493_));
  NOR4_X1   g292(.A1(new_n482_), .A2(new_n474_), .A3(KEYINPUT33), .A4(new_n479_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n488_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n433_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n395_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n469_), .A2(new_n470_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n473_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n471_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n473_), .A2(new_n500_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n499_), .B(new_n479_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n487_), .A2(new_n396_), .A3(new_n488_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n498_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  OAI22_X1  g305(.A1(new_n441_), .A2(new_n490_), .B1(new_n495_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT87), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G228gat), .A2(G233gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT84), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n464_), .A2(KEYINPUT29), .B1(new_n508_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n410_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n511_), .A2(new_n508_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n410_), .A2(new_n512_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G78gat), .B(G106gat), .Z(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n515_), .A2(new_n521_), .A3(new_n517_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n464_), .A2(KEYINPUT29), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT28), .B(G22gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G50gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n523_), .B(new_n525_), .ZN(new_n526_));
  AND4_X1   g325(.A1(KEYINPUT88), .A2(new_n520_), .A3(new_n522_), .A4(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT88), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n529_), .A2(new_n526_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n507_), .A2(new_n532_), .A3(KEYINPUT93), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n395_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(KEYINPUT27), .A3(new_n505_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n484_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n498_), .A2(new_n505_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT27), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n531_), .A2(new_n535_), .A3(new_n536_), .A4(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT93), .B1(new_n507_), .B2(new_n532_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n391_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n535_), .A2(new_n539_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n531_), .A2(new_n391_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n544_), .A2(new_n536_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT94), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n271_), .A2(new_n238_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n241_), .B2(new_n271_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT75), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n271_), .B(new_n238_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n551_), .A2(new_n552_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n553_), .B1(new_n560_), .B2(KEYINPUT75), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G169gat), .B(G197gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n561_), .B(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n548_), .A2(new_n549_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n498_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n481_), .A2(KEYINPUT33), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n492_), .A2(new_n491_), .A3(new_n480_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n496_), .A2(new_n497_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n573_), .A2(new_n397_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT32), .B(new_n396_), .C1(new_n435_), .C2(new_n439_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n569_), .A2(new_n572_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n568_), .B1(new_n576_), .B2(new_n531_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(new_n533_), .A3(new_n540_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n546_), .B1(new_n578_), .B2(new_n391_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n566_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT94), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  AOI211_X1 g380(.A(new_n299_), .B(new_n336_), .C1(new_n567_), .C2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(new_n266_), .A3(new_n484_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT38), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n582_), .A2(new_n266_), .A3(new_n484_), .A4(new_n585_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n263_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT97), .B1(new_n548_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT97), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n579_), .A2(new_n591_), .A3(new_n263_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n335_), .A2(new_n566_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(new_n297_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n593_), .A2(new_n536_), .A3(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n587_), .B(new_n588_), .C1(new_n597_), .C2(new_n266_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT98), .ZN(G1324gat));
  INV_X1    g398(.A(new_n544_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n582_), .A2(new_n267_), .A3(new_n600_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n600_), .B(new_n595_), .C1(new_n590_), .C2(new_n592_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n267_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n605_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n601_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT40), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(KEYINPUT40), .B(new_n601_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1325gat));
  INV_X1    g412(.A(G15gat), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n593_), .A2(new_n596_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n391_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT41), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n582_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(G1326gat));
  INV_X1    g421(.A(G22gat), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n615_), .B2(new_n531_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT42), .Z(new_n625_));
  NAND3_X1  g424(.A1(new_n582_), .A2(new_n623_), .A3(new_n531_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1327gat));
  INV_X1    g426(.A(new_n297_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n589_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI211_X1 g429(.A(new_n336_), .B(new_n630_), .C1(new_n567_), .C2(new_n581_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n632_), .A2(G29gat), .A3(new_n536_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n594_), .A2(new_n628_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n548_), .B2(new_n264_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n264_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n579_), .A2(KEYINPUT43), .A3(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT44), .B(new_n634_), .C1(new_n636_), .C2(new_n638_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n484_), .A3(new_n642_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(KEYINPUT100), .A3(G29gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT100), .B1(new_n643_), .B2(G29gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n633_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT101), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n633_), .B(new_n648_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1328gat));
  NOR2_X1   g449(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n641_), .A2(new_n600_), .A3(new_n642_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n641_), .A2(KEYINPUT102), .A3(new_n600_), .A4(new_n642_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n654_), .A2(G36gat), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT45), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n544_), .A2(G36gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n631_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n567_), .A2(new_n581_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n661_), .A2(new_n335_), .A3(new_n629_), .A4(new_n659_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(KEYINPUT103), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n657_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n631_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(KEYINPUT103), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(KEYINPUT45), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n651_), .B1(new_n656_), .B2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n654_), .A2(G36gat), .A3(new_n655_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n651_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n670_), .A2(new_n671_), .A3(new_n667_), .A4(new_n664_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n672_), .ZN(G1329gat));
  NOR3_X1   g472(.A1(new_n632_), .A2(G43gat), .A3(new_n391_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n641_), .A2(new_n616_), .A3(new_n642_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(G43gat), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g476(.A1(new_n632_), .A2(G50gat), .A3(new_n532_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n641_), .A2(new_n531_), .A3(new_n642_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n680_), .A3(G50gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n679_), .B2(G50gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT106), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n678_), .B(new_n685_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1331gat));
  NOR2_X1   g486(.A1(new_n335_), .A2(new_n566_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n548_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n299_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n484_), .ZN(new_n691_));
  NOR4_X1   g490(.A1(new_n593_), .A2(new_n297_), .A3(new_n335_), .A4(new_n566_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n274_), .B1(new_n484_), .B2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n693_), .B2(new_n274_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n691_), .B1(new_n692_), .B2(new_n695_), .ZN(G1332gat));
  AOI21_X1  g495(.A(new_n275_), .B1(new_n692_), .B2(new_n600_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT48), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n690_), .A2(new_n275_), .A3(new_n600_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1333gat));
  INV_X1    g499(.A(G71gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n692_), .B2(new_n616_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT49), .Z(new_n703_));
  NAND2_X1  g502(.A1(new_n616_), .A2(new_n701_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT108), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n690_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1334gat));
  INV_X1    g506(.A(G78gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n692_), .B2(new_n531_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT50), .Z(new_n710_));
  NAND3_X1  g509(.A1(new_n690_), .A2(new_n708_), .A3(new_n531_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1335gat));
  NAND3_X1  g511(.A1(new_n548_), .A2(new_n629_), .A3(new_n688_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n484_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n636_), .A2(new_n638_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n688_), .A2(new_n297_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n536_), .A2(new_n217_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(G1336gat));
  AOI21_X1  g519(.A(G92gat), .B1(new_n714_), .B2(new_n600_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n544_), .A2(new_n218_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n718_), .B2(new_n722_), .ZN(G1337gat));
  NAND3_X1  g522(.A1(new_n714_), .A2(new_n214_), .A3(new_n616_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n718_), .A2(new_n616_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(G99gat), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT109), .B(new_n227_), .C1(new_n718_), .C2(new_n616_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT51), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n731_), .B(new_n724_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1338gat));
  NAND3_X1  g532(.A1(new_n714_), .A2(new_n215_), .A3(new_n531_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n718_), .A2(new_n531_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G106gat), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT52), .B(new_n228_), .C1(new_n718_), .C2(new_n531_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT111), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n734_), .B(new_n741_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1339gat));
  NAND3_X1  g544(.A1(new_n298_), .A2(new_n335_), .A3(new_n580_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT54), .Z(new_n747_));
  AND2_X1   g546(.A1(new_n566_), .A2(new_n332_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n309_), .A2(new_n753_), .A3(new_n318_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n308_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(KEYINPUT112), .A2(G230gat), .A3(G233gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n756_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n308_), .A2(new_n315_), .A3(new_n316_), .A4(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n307_), .A2(new_n753_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n754_), .A2(KEYINPUT113), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n330_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT113), .B1(new_n754_), .B2(new_n761_), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT114), .B(new_n752_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n763_), .A2(new_n750_), .A3(new_n764_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(KEYINPUT115), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n754_), .A2(new_n761_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(new_n330_), .A3(new_n762_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n752_), .B1(new_n771_), .B2(KEYINPUT114), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n748_), .B1(new_n767_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n331_), .A2(new_n332_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n556_), .A2(new_n552_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n565_), .B1(new_n551_), .B2(new_n557_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n561_), .A2(new_n565_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n773_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n589_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n778_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT114), .B1(new_n763_), .B2(new_n764_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n751_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n770_), .A2(KEYINPUT56), .A3(new_n330_), .A4(new_n762_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n749_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n784_), .A2(new_n786_), .A3(new_n765_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n782_), .B1(new_n787_), .B2(new_n748_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT116), .B1(new_n788_), .B2(new_n263_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n781_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n263_), .B1(new_n773_), .B2(new_n778_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT57), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n777_), .A2(new_n332_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n750_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n797_));
  AOI211_X1 g596(.A(new_n795_), .B(new_n796_), .C1(new_n797_), .C2(new_n785_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n785_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n264_), .B1(new_n799_), .B2(KEYINPUT58), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n800_), .B2(KEYINPUT117), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n264_), .B(new_n802_), .C1(new_n799_), .C2(KEYINPUT58), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n794_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(KEYINPUT117), .ZN(new_n805_));
  INV_X1    g604(.A(new_n798_), .ZN(new_n806_));
  AND4_X1   g605(.A1(new_n794_), .A2(new_n805_), .A3(new_n803_), .A4(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n791_), .B(new_n793_), .C1(new_n804_), .C2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n747_), .B1(new_n808_), .B2(new_n297_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n544_), .A2(new_n545_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(new_n536_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT59), .B1(new_n809_), .B2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(KEYINPUT59), .ZN(new_n815_));
  INV_X1    g614(.A(new_n747_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(KEYINPUT57), .A2(new_n792_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n628_), .B1(new_n791_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n816_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT119), .B(new_n628_), .C1(new_n791_), .C2(new_n817_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n815_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n566_), .A2(G113gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT120), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n814_), .A2(new_n822_), .A3(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n790_), .B1(new_n792_), .B2(new_n780_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n788_), .A2(KEYINPUT116), .A3(new_n263_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n793_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n807_), .A2(new_n804_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n297_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n816_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n566_), .A3(new_n812_), .ZN(new_n832_));
  INV_X1    g631(.A(G113gat), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n825_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n825_), .A2(new_n834_), .A3(KEYINPUT121), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(G1340gat));
  NAND3_X1  g638(.A1(new_n814_), .A2(new_n822_), .A3(new_n336_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G120gat), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n809_), .A2(new_n813_), .ZN(new_n842_));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n335_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n842_), .B(new_n844_), .C1(KEYINPUT60), .C2(new_n843_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n845_), .ZN(G1341gat));
  NAND4_X1  g645(.A1(new_n747_), .A2(new_n628_), .A3(new_n484_), .A4(new_n810_), .ZN(new_n847_));
  INV_X1    g646(.A(G127gat), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n847_), .A2(KEYINPUT122), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT122), .B1(new_n847_), .B2(new_n848_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n814_), .A2(new_n822_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n297_), .A2(new_n848_), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n849_), .B(new_n850_), .C1(new_n851_), .C2(new_n852_), .ZN(G1342gat));
  AOI21_X1  g652(.A(G134gat), .B1(new_n842_), .B2(new_n263_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n264_), .A2(G134gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT123), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n851_), .B2(new_n856_), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n532_), .A2(new_n616_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n831_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n600_), .A2(new_n536_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n859_), .A2(new_n580_), .A3(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n447_), .ZN(G1344gat));
  NOR3_X1   g662(.A1(new_n859_), .A2(new_n335_), .A3(new_n861_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(new_n448_), .ZN(G1345gat));
  NAND4_X1  g664(.A1(new_n831_), .A2(new_n628_), .A3(new_n858_), .A4(new_n860_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT124), .ZN(new_n867_));
  INV_X1    g666(.A(new_n858_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n830_), .B2(new_n816_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT124), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n628_), .A4(new_n860_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n867_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n867_), .B2(new_n871_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1346gat));
  NOR2_X1   g674(.A1(new_n859_), .A2(new_n861_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G162gat), .B1(new_n876_), .B2(new_n263_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n264_), .A2(G162gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n876_), .B2(new_n878_), .ZN(G1347gat));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n544_), .A2(new_n484_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n391_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n531_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n566_), .B(new_n885_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n880_), .B1(new_n887_), .B2(new_n340_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n886_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n338_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(G1348gat));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n336_), .B(new_n885_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n894_), .B2(G176gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n893_), .A2(KEYINPUT125), .A3(new_n342_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n809_), .A2(new_n531_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n884_), .A2(new_n335_), .A3(new_n342_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n895_), .A2(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(G1349gat));
  OR2_X1    g698(.A1(new_n820_), .A2(new_n821_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n900_), .A2(new_n885_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n297_), .B1(new_n360_), .B2(new_n418_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n897_), .A2(new_n628_), .A3(new_n883_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n901_), .A2(new_n902_), .B1(new_n903_), .B2(new_n348_), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n901_), .A2(new_n263_), .A3(new_n417_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n264_), .B(new_n885_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(G190gat), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n907_), .A2(new_n906_), .A3(G190gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n905_), .B1(new_n908_), .B2(new_n909_), .ZN(G1351gat));
  NAND3_X1  g709(.A1(new_n869_), .A2(new_n566_), .A3(new_n881_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g711(.A1(new_n859_), .A2(new_n335_), .A3(new_n882_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(KEYINPUT127), .B2(new_n326_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT127), .B(G204gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n913_), .B2(new_n915_), .ZN(G1353gat));
  NAND3_X1  g715(.A1(new_n869_), .A2(new_n628_), .A3(new_n881_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AND2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n920_), .B1(new_n917_), .B2(new_n918_), .ZN(G1354gat));
  NOR2_X1   g720(.A1(new_n859_), .A2(new_n882_), .ZN(new_n922_));
  AOI21_X1  g721(.A(G218gat), .B1(new_n922_), .B2(new_n263_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n264_), .A2(G218gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(new_n924_), .ZN(G1355gat));
endmodule


