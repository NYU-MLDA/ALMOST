//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_, new_n966_;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G92gat), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT9), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n208_), .A2(new_n211_), .A3(new_n216_), .A4(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n209_), .A2(new_n210_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n214_), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n218_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n224_), .B1(new_n227_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT8), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n231_), .B(new_n230_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n224_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n222_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G57gat), .B(G64gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G78gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(KEYINPUT11), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n242_));
  INV_X1    g041(.A(new_n240_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n241_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n238_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n231_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AOI211_X1 g049(.A(KEYINPUT8), .B(new_n223_), .C1(new_n250_), .C2(new_n216_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n236_), .B1(new_n235_), .B2(new_n224_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n246_), .B(new_n221_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n204_), .B1(new_n247_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT65), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n221_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT66), .B(new_n221_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n260_));
  OAI211_X1 g059(.A(KEYINPUT12), .B(new_n241_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n259_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT12), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(new_n238_), .B2(new_n246_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n263_), .A2(new_n203_), .A3(new_n253_), .A4(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n246_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n257_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n253_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n204_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G120gat), .B(G148gat), .Z(new_n272_));
  XNOR2_X1  g071(.A(G176gat), .B(G204gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n256_), .A2(new_n266_), .A3(new_n271_), .A4(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n270_), .B1(new_n269_), .B2(new_n204_), .ZN(new_n280_));
  AOI211_X1 g079(.A(KEYINPUT65), .B(new_n203_), .C1(new_n268_), .C2(new_n253_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n282_), .A2(KEYINPUT68), .A3(new_n266_), .A4(new_n276_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n266_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n276_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(KEYINPUT13), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT13), .B1(new_n284_), .B2(new_n287_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n202_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n287_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT13), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(KEYINPUT69), .A3(new_n288_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(G197gat), .A2(G204gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G197gat), .A2(G204gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(KEYINPUT90), .A2(KEYINPUT21), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(KEYINPUT89), .A2(G211gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(KEYINPUT89), .A2(G211gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(G218gat), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(KEYINPUT89), .A2(G211gat), .ZN(new_n305_));
  INV_X1    g104(.A(G218gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(KEYINPUT89), .A2(G211gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n301_), .A2(new_n304_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n301_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n298_), .A2(new_n299_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n308_), .B(new_n304_), .C1(new_n312_), .C2(KEYINPUT21), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n310_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT3), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT86), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT87), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n315_), .A2(KEYINPUT86), .A3(new_n316_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n321_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT85), .B1(new_n333_), .B2(KEYINPUT1), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT85), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(G155gat), .A4(G162gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n333_), .A2(KEYINPUT1), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n336_), .A2(new_n339_), .A3(new_n340_), .A4(new_n332_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n315_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n342_), .A2(new_n322_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n331_), .A2(new_n335_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n314_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G228gat), .ZN(new_n347_));
  OR2_X1    g146(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G78gat), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n351_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n218_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(G106gat), .A3(new_n353_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n346_), .B(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n318_), .A2(new_n319_), .ZN(new_n359_));
  INV_X1    g158(.A(G141gat), .ZN(new_n360_));
  INV_X1    g159(.A(G148gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n316_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n364_), .A3(new_n330_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n327_), .B(new_n325_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n335_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n341_), .A2(new_n343_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT28), .B1(new_n369_), .B2(KEYINPUT29), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n344_), .A2(new_n371_), .A3(new_n345_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G22gat), .B(G50gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n371_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n376_));
  AND4_X1   g175(.A1(new_n371_), .A2(new_n367_), .A3(new_n345_), .A4(new_n368_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n358_), .A2(KEYINPUT91), .A3(new_n374_), .A4(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(KEYINPUT91), .A3(new_n374_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n313_), .A2(new_n311_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n309_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n369_), .B2(KEYINPUT29), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(new_n357_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT91), .B1(new_n378_), .B2(new_n374_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n379_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G183gat), .ZN(new_n388_));
  INV_X1    g187(.A(G190gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT23), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(G183gat), .A3(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(G183gat), .B2(G190gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G169gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n391_), .B1(G183gat), .B2(G190gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(KEYINPUT82), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n400_), .A2(new_n391_), .A3(G183gat), .A4(G190gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n398_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G169gat), .ZN(new_n403_));
  INV_X1    g202(.A(G176gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(KEYINPUT80), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(G169gat), .B2(G176gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT24), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n402_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT24), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(G169gat), .B2(G176gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT26), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(G190gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT78), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n388_), .A3(KEYINPUT25), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n389_), .A2(KEYINPUT79), .A3(KEYINPUT26), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT25), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT78), .B1(new_n420_), .B2(G183gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(G183gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n414_), .A2(G190gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(KEYINPUT81), .B(new_n412_), .C1(new_n419_), .C2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n409_), .A2(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n427_));
  OAI22_X1  g226(.A1(KEYINPUT25), .A2(new_n388_), .B1(new_n389_), .B2(KEYINPUT26), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n416_), .B1(KEYINPUT25), .B2(new_n388_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT81), .B1(new_n431_), .B2(new_n412_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n397_), .B1(new_n426_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n314_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G183gat), .A2(G190gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n396_), .B1(new_n402_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n408_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT25), .B(G183gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT26), .B(G190gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n437_), .A2(new_n440_), .A3(new_n393_), .A4(new_n412_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT92), .B1(new_n314_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT92), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n382_), .A2(new_n444_), .A3(new_n436_), .A4(new_n441_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT19), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n434_), .A2(new_n443_), .A3(new_n445_), .A4(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n314_), .B2(new_n442_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n382_), .B(new_n397_), .C1(new_n426_), .C2(new_n432_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n447_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G8gat), .B(G36gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(G64gat), .B(G92gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT32), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n450_), .A2(new_n454_), .A3(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G127gat), .B(G134gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G113gat), .B(G120gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR4_X1   g264(.A1(new_n363_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n466_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n334_), .B1(new_n467_), .B2(new_n329_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n368_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n465_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n367_), .A2(new_n368_), .A3(new_n464_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(KEYINPUT4), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G225gat), .A2(G233gat), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n464_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT4), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n470_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G29gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G85gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT0), .B(G57gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n477_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n461_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT97), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n412_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT81), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n425_), .A3(new_n409_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n382_), .B1(new_n491_), .B2(new_n397_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n314_), .B2(new_n442_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n447_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n447_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n451_), .A2(new_n452_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n460_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n487_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI211_X1 g301(.A(KEYINPUT97), .B(new_n460_), .C1(new_n496_), .C2(new_n498_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n486_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n473_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n470_), .A2(new_n471_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n482_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT95), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(KEYINPUT95), .A3(new_n482_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n506_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n472_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n367_), .A2(new_n368_), .A3(new_n464_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n515_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n506_), .B1(new_n470_), .B2(KEYINPUT4), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n478_), .B(new_n483_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n477_), .A2(new_n478_), .A3(new_n483_), .A4(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n514_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n459_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n445_), .A2(new_n449_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n436_), .A2(new_n441_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n444_), .B1(new_n526_), .B2(new_n382_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n525_), .A2(new_n527_), .A3(new_n492_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n497_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n524_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n450_), .A2(new_n454_), .A3(new_n459_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n523_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n387_), .B1(new_n505_), .B2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n380_), .A2(new_n384_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n380_), .A2(new_n384_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n386_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT27), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n450_), .A2(new_n454_), .A3(new_n459_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n459_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n477_), .A2(new_n478_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n482_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n518_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n499_), .A2(new_n524_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(KEYINPUT27), .A3(new_n531_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n538_), .A2(new_n542_), .A3(new_n546_), .A4(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n534_), .A2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT84), .B(G43gat), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n491_), .A2(new_n397_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(new_n491_), .B2(new_n397_), .ZN(new_n554_));
  INV_X1    g353(.A(G71gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G227gat), .A2(G233gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(G15gat), .ZN(new_n557_));
  INV_X1    g356(.A(G15gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(G227gat), .A3(G233gat), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n555_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(new_n559_), .A3(new_n555_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(G99gat), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n229_), .B1(new_n564_), .B2(new_n560_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n563_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n569_));
  OAI22_X1  g368(.A1(new_n553_), .A2(new_n554_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n433_), .A2(new_n551_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n491_), .A2(new_n397_), .A3(new_n552_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n568_), .A2(new_n569_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n570_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n571_), .B1(new_n570_), .B2(new_n575_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n464_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n574_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT31), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n570_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n465_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n546_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n542_), .A2(new_n387_), .A3(new_n548_), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT98), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n464_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n581_), .A2(new_n465_), .A3(new_n582_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n545_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n525_), .A2(new_n527_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n529_), .B1(new_n591_), .B2(new_n434_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n539_), .B1(new_n592_), .B2(new_n459_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n539_), .A2(new_n532_), .B1(new_n593_), .B2(new_n547_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n590_), .A2(new_n594_), .A3(new_n595_), .A4(new_n387_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n550_), .A2(new_n584_), .B1(new_n587_), .B2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G15gat), .B(G22gat), .ZN(new_n598_));
  INV_X1    g397(.A(G1gat), .ZN(new_n599_));
  INV_X1    g398(.A(G8gat), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT14), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G1gat), .B(G8gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G29gat), .B(G36gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G43gat), .B(G50gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n604_), .B(new_n607_), .Z(new_n608_));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n607_), .B(KEYINPUT15), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(new_n604_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n604_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n607_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n609_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n611_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT77), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G113gat), .B(G141gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G169gat), .B(G197gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n620_), .B(new_n621_), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n619_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(KEYINPUT36), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n238_), .A2(new_n607_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT71), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n631_));
  NAND2_X1  g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n631_), .B(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n634_), .B2(KEYINPUT35), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n631_), .B(new_n632_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT35), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(KEYINPUT71), .A3(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  AOI22_X1  g438(.A1(new_n635_), .A2(new_n638_), .B1(new_n639_), .B2(KEYINPUT72), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n629_), .A2(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n639_), .A2(KEYINPUT72), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n259_), .A2(new_n612_), .A3(new_n260_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n641_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n642_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n628_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n646_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n627_), .B(KEYINPUT36), .Z(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n644_), .A3(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n650_), .A3(KEYINPUT37), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT73), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n653_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n648_), .A2(KEYINPUT73), .A3(new_n644_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n649_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n647_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT37), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n652_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(G127gat), .B(G155gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT16), .ZN(new_n661_));
  XNOR2_X1  g460(.A(G183gat), .B(G211gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT17), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT75), .Z(new_n665_));
  NAND2_X1  g464(.A1(G231gat), .A2(G233gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n604_), .B(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(new_n267_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT74), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n667_), .B(new_n246_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(KEYINPUT74), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n665_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n663_), .B(KEYINPUT17), .Z(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT76), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT76), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n671_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n673_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n659_), .A2(new_n679_), .ZN(new_n680_));
  NOR4_X1   g479(.A1(new_n297_), .A2(new_n597_), .A3(new_n624_), .A4(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n599_), .A3(new_n545_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT38), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT99), .Z(new_n685_));
  INV_X1    g484(.A(new_n657_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n597_), .A2(new_n686_), .ZN(new_n687_));
  AND4_X1   g486(.A1(new_n623_), .A2(new_n687_), .A3(new_n296_), .A4(new_n679_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n599_), .B1(new_n688_), .B2(new_n545_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n683_), .B2(new_n682_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n685_), .A2(new_n690_), .ZN(G1324gat));
  INV_X1    g490(.A(new_n594_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G8gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT39), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n681_), .A2(new_n600_), .A3(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1325gat));
  INV_X1    g498(.A(new_n584_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n558_), .B1(new_n688_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT41), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n681_), .A2(new_n558_), .A3(new_n700_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1326gat));
  INV_X1    g503(.A(G22gat), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n538_), .B(KEYINPUT101), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n688_), .B2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT42), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n681_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1327gat));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n686_), .A2(new_n678_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT105), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(new_n296_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n597_), .A2(new_n624_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n716_), .A2(G29gat), .A3(new_n546_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n289_), .A2(new_n290_), .A3(new_n202_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT69), .B1(new_n294_), .B2(new_n288_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n623_), .B(new_n678_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n296_), .A2(KEYINPUT102), .A3(new_n623_), .A4(new_n678_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n597_), .B2(new_n659_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n587_), .A2(new_n596_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n540_), .A2(new_n541_), .ZN(new_n728_));
  AOI22_X1  g527(.A1(new_n508_), .A2(new_n509_), .B1(new_n472_), .B2(new_n512_), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n484_), .A2(new_n521_), .B1(new_n729_), .B2(new_n511_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n728_), .A2(new_n730_), .A3(new_n520_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n545_), .B(new_n461_), .C1(new_n501_), .C2(new_n503_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n538_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  AND4_X1   g532(.A1(new_n538_), .A2(new_n546_), .A3(new_n542_), .A4(new_n548_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n584_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT43), .B(new_n659_), .C1(new_n727_), .C2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n726_), .B1(new_n736_), .B2(KEYINPUT103), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n727_), .A2(new_n735_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n739_));
  INV_X1    g538(.A(new_n659_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n725_), .B(KEYINPUT44), .C1(new_n737_), .C2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n725_), .B1(new_n737_), .B2(new_n743_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT44), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n736_), .A2(KEYINPUT103), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n741_), .A2(new_n742_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n726_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(KEYINPUT104), .A3(new_n725_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n745_), .B1(new_n748_), .B2(new_n752_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(new_n545_), .ZN(new_n754_));
  INV_X1    g553(.A(G29gat), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n711_), .B(new_n718_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n753_), .B2(new_n545_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT106), .B1(new_n757_), .B2(new_n717_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1328gat));
  INV_X1    g558(.A(new_n716_), .ZN(new_n760_));
  INV_X1    g559(.A(G36gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n692_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT45), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n753_), .A2(new_n692_), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT46), .B(new_n763_), .C1(new_n764_), .C2(new_n761_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n766_));
  INV_X1    g565(.A(new_n763_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n761_), .B1(new_n753_), .B2(new_n692_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n769_), .ZN(G1329gat));
  AOI21_X1  g569(.A(G43gat), .B1(new_n760_), .B2(new_n700_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT108), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n746_), .A2(new_n747_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n752_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n700_), .A2(G43gat), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n744_), .A2(new_n776_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n775_), .A2(KEYINPUT107), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT107), .B1(new_n775_), .B2(new_n777_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n772_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT47), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n772_), .B(new_n782_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1330gat));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n753_), .A2(new_n785_), .A3(new_n538_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(G50gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n753_), .B2(new_n538_), .ZN(new_n788_));
  INV_X1    g587(.A(G50gat), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n706_), .A2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT110), .ZN(new_n791_));
  OAI22_X1  g590(.A1(new_n787_), .A2(new_n788_), .B1(new_n716_), .B2(new_n791_), .ZN(G1331gat));
  NOR2_X1   g591(.A1(new_n597_), .A2(new_n623_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n296_), .A2(new_n680_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(KEYINPUT111), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(KEYINPUT111), .B2(new_n794_), .ZN(new_n796_));
  INV_X1    g595(.A(G57gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n545_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n679_), .A2(new_n624_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n296_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n687_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G57gat), .B1(new_n801_), .B2(new_n546_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n798_), .A2(new_n802_), .ZN(G1332gat));
  OAI21_X1  g602(.A(G64gat), .B1(new_n801_), .B2(new_n594_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT48), .ZN(new_n805_));
  INV_X1    g604(.A(G64gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n796_), .A2(new_n806_), .A3(new_n692_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1333gat));
  OAI21_X1  g607(.A(G71gat), .B1(new_n801_), .B2(new_n584_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT49), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n796_), .A2(new_n555_), .A3(new_n700_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1334gat));
  NAND3_X1  g611(.A1(new_n796_), .A2(new_n351_), .A3(new_n706_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n800_), .A2(new_n687_), .A3(new_n706_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(G78gat), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT50), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(G1335gat));
  AND3_X1   g616(.A1(new_n793_), .A2(new_n297_), .A3(new_n713_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n206_), .A3(new_n545_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n296_), .A2(new_n623_), .A3(new_n679_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n751_), .A2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT112), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n822_), .A2(new_n545_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n819_), .B1(new_n823_), .B2(new_n206_), .ZN(G1336gat));
  AOI21_X1  g623(.A(G92gat), .B1(new_n818_), .B2(new_n692_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n692_), .A2(new_n205_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT113), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n822_), .B2(new_n827_), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT114), .Z(G1337gat));
  NAND3_X1  g628(.A1(new_n751_), .A2(new_n700_), .A3(new_n820_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n700_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n830_), .A2(G99gat), .B1(new_n818_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(KEYINPUT115), .B2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(KEYINPUT115), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(G1338gat));
  NAND3_X1  g635(.A1(new_n818_), .A2(new_n218_), .A3(new_n538_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n751_), .A2(new_n538_), .A3(new_n820_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(KEYINPUT117), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n218_), .B1(new_n839_), .B2(KEYINPUT117), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n838_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n838_), .B2(new_n841_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n837_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g644(.A1(new_n692_), .A2(new_n546_), .A3(new_n584_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n617_), .A2(new_n622_), .ZN(new_n847_));
  AOI211_X1 g646(.A(new_n609_), .B(new_n613_), .C1(new_n614_), .C2(new_n607_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n849_), .B2(new_n622_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n254_), .B1(new_n264_), .B2(new_n268_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n203_), .B1(new_n851_), .B2(new_n263_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n266_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n851_), .A2(KEYINPUT55), .A3(new_n203_), .A4(new_n263_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n856_), .A2(KEYINPUT56), .A3(new_n286_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT56), .B1(new_n856_), .B2(new_n286_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n284_), .B(new_n850_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861_));
  OR3_X1    g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n659_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n292_), .A2(new_n850_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n284_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n624_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n657_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n868_), .A2(KEYINPUT57), .A3(new_n657_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n865_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n873_), .A2(new_n678_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n799_), .B(KEYINPUT118), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n289_), .A2(new_n290_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT54), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n875_), .A2(new_n876_), .A3(new_n659_), .A4(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n877_), .A2(KEYINPUT54), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n387_), .B(new_n846_), .C1(new_n874_), .C2(new_n881_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n880_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n879_), .B(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n873_), .A2(new_n678_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(KEYINPUT121), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n888_), .A2(new_n387_), .A3(new_n846_), .A4(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n884_), .A2(new_n623_), .A3(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G113gat), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n624_), .A2(G113gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n882_), .B2(new_n895_), .ZN(G1340gat));
  NAND3_X1  g695(.A1(new_n884_), .A2(new_n297_), .A3(new_n892_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G120gat), .ZN(new_n898_));
  INV_X1    g697(.A(new_n888_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n538_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n901_));
  AOI21_X1  g700(.A(G120gat), .B1(new_n297_), .B2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n901_), .B2(G120gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n900_), .A2(new_n846_), .A3(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n898_), .A2(new_n904_), .ZN(G1341gat));
  INV_X1    g704(.A(G127gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n678_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n884_), .A2(new_n892_), .A3(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n882_), .B2(new_n678_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n908_), .A2(KEYINPUT122), .A3(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(KEYINPUT122), .B1(new_n908_), .B2(new_n909_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1342gat));
  XNOR2_X1  g711(.A(KEYINPUT123), .B(G134gat), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n884_), .A2(new_n740_), .A3(new_n892_), .A4(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(G134gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n915_), .B1(new_n882_), .B2(new_n657_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1343gat));
  NAND4_X1  g716(.A1(new_n584_), .A2(new_n594_), .A3(new_n538_), .A4(new_n545_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n899_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n623_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n297_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g722(.A1(new_n919_), .A2(new_n679_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT61), .B(G155gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1346gat));
  INV_X1    g725(.A(G162gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n919_), .A2(new_n927_), .A3(new_n686_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n899_), .A2(new_n659_), .A3(new_n918_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(G1347gat));
  XNOR2_X1  g729(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n706_), .A2(new_n594_), .A3(new_n585_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n888_), .A2(new_n623_), .A3(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n933_), .B2(KEYINPUT22), .ZN(new_n934_));
  OAI21_X1  g733(.A(G169gat), .B1(new_n933_), .B2(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n403_), .B2(new_n934_), .ZN(G1348gat));
  AND2_X1   g736(.A1(new_n888_), .A2(new_n932_), .ZN(new_n938_));
  AOI21_X1  g737(.A(G176gat), .B1(new_n938_), .B2(new_n297_), .ZN(new_n939_));
  NOR4_X1   g738(.A1(new_n296_), .A2(new_n404_), .A3(new_n594_), .A4(new_n585_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(new_n900_), .B2(new_n940_), .ZN(G1349gat));
  NAND4_X1  g740(.A1(new_n900_), .A2(new_n692_), .A3(new_n590_), .A4(new_n679_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n678_), .A2(new_n438_), .ZN(new_n943_));
  AOI22_X1  g742(.A1(new_n942_), .A2(new_n388_), .B1(new_n938_), .B2(new_n943_), .ZN(G1350gat));
  NAND2_X1  g743(.A1(new_n686_), .A2(new_n439_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(KEYINPUT125), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n938_), .A2(new_n946_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n938_), .A2(new_n740_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n389_), .ZN(G1351gat));
  NAND4_X1  g748(.A1(new_n692_), .A2(new_n538_), .A3(new_n546_), .A4(new_n584_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n899_), .A2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(new_n623_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(G204gat), .ZN(new_n955_));
  XOR2_X1   g754(.A(KEYINPUT126), .B(G204gat), .Z(new_n956_));
  NAND2_X1  g755(.A1(new_n951_), .A2(new_n297_), .ZN(new_n957_));
  MUX2_X1   g756(.A(new_n955_), .B(new_n956_), .S(new_n957_), .Z(G1353gat));
  NAND2_X1  g757(.A1(new_n951_), .A2(new_n679_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  AND2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n959_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n962_), .B1(new_n959_), .B2(new_n960_), .ZN(G1354gat));
  AOI21_X1  g762(.A(G218gat), .B1(new_n951_), .B2(new_n686_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n659_), .A2(new_n306_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(KEYINPUT127), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n964_), .B1(new_n951_), .B2(new_n966_), .ZN(G1355gat));
endmodule


