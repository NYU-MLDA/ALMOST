//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209_));
  XNOR2_X1  g008(.A(G29gat), .B(G36gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n213_), .B(KEYINPUT15), .Z(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(new_n208_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n208_), .B(new_n213_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n217_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n218_), .B1(KEYINPUT77), .B2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n222_), .B1(KEYINPUT77), .B2(new_n221_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT78), .B(G113gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(G141gat), .ZN(new_n225_));
  XOR2_X1   g024(.A(G169gat), .B(G197gat), .Z(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n223_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230_));
  INV_X1    g029(.A(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT7), .ZN(new_n234_));
  AND3_X1   g033(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n230_), .A2(new_n238_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n234_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n241_));
  INV_X1    g040(.A(G85gat), .ZN(new_n242_));
  INV_X1    g041(.A(G92gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G85gat), .A2(G92gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n240_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT8), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n241_), .B1(new_n240_), .B2(new_n246_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(new_n246_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT8), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(KEYINPUT65), .A3(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n244_), .A2(KEYINPUT9), .A3(new_n245_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n245_), .A2(KEYINPUT9), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n237_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT10), .B(G99gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(G106gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n253_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT66), .B1(new_n250_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n251_), .A2(KEYINPUT65), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(KEYINPUT8), .A3(new_n247_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n259_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G71gat), .B(G78gat), .Z(new_n269_));
  INV_X1    g068(.A(G57gat), .ZN(new_n270_));
  INV_X1    g069(.A(G64gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G57gat), .A2(G64gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT11), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT67), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n281_), .A3(KEYINPUT11), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n277_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n268_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n262_), .A2(new_n288_), .A3(new_n267_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(G230gat), .A3(G233gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT12), .B1(new_n284_), .B2(new_n285_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(new_n266_), .B2(new_n264_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n268_), .B2(new_n286_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G230gat), .A2(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT12), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n289_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n291_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G176gat), .B(G204gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(G120gat), .B(G148gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n299_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n291_), .A2(new_n298_), .A3(new_n304_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT13), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n306_), .B(new_n307_), .C1(KEYINPUT69), .C2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G190gat), .B(G218gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G134gat), .B(G162gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  INV_X1    g116(.A(KEYINPUT36), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G232gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT34), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n321_), .A2(KEYINPUT35), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n213_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n264_), .A2(new_n266_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n215_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n322_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n213_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n265_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n215_), .A2(new_n324_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n321_), .A2(KEYINPUT35), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n322_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n330_), .A2(KEYINPUT70), .A3(new_n331_), .A4(new_n333_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n319_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT37), .B1(new_n338_), .B2(KEYINPUT72), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n317_), .B(KEYINPUT36), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n341_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n336_), .A2(new_n337_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n337_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n330_), .A2(new_n331_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT70), .B1(new_n346_), .B2(new_n322_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n347_), .B2(new_n334_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n344_), .B1(new_n348_), .B2(new_n319_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n339_), .B(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G231gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n208_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(new_n286_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT74), .ZN(new_n354_));
  XOR2_X1   g153(.A(G183gat), .B(G211gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(G127gat), .B(G155gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT17), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT75), .Z(new_n362_));
  INV_X1    g161(.A(KEYINPUT17), .ZN(new_n363_));
  OR3_X1    g162(.A1(new_n353_), .A2(new_n363_), .A3(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n314_), .A2(new_n350_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n229_), .B1(new_n366_), .B2(KEYINPUT76), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT30), .B(G99gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373_));
  NAND3_X1  g172(.A1(KEYINPUT80), .A2(G183gat), .A3(G190gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n378_));
  NAND2_X1  g177(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n370_), .A3(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n372_), .A2(KEYINPUT81), .A3(new_n373_), .A4(new_n374_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT24), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385_));
  MUX2_X1   g184(.A(new_n384_), .B(KEYINPUT24), .S(new_n385_), .Z(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT26), .B(G190gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n387_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n382_), .A2(new_n386_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G176gat), .ZN(new_n393_));
  AND2_X1   g192(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n396_), .A2(new_n383_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n373_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n370_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n378_), .A2(new_n379_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G183gat), .A2(G190gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n397_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n369_), .B1(new_n392_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  INV_X1    g205(.A(G71gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n392_), .A2(new_n403_), .A3(new_n369_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n410_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n408_), .B1(new_n412_), .B2(new_n404_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n368_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n414_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n409_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n412_), .A2(new_n408_), .A3(new_n404_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(KEYINPUT84), .A3(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(KEYINPUT82), .A2(KEYINPUT83), .ZN(new_n424_));
  NAND2_X1  g223(.A1(KEYINPUT82), .A2(KEYINPUT83), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G127gat), .A2(G134gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G127gat), .A2(G134gat), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n424_), .B(new_n425_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(G127gat), .A2(G134gat), .ZN(new_n430_));
  AND2_X1   g229(.A1(KEYINPUT82), .A2(KEYINPUT83), .ZN(new_n431_));
  NOR2_X1   g230(.A1(KEYINPUT82), .A2(KEYINPUT83), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n430_), .B(new_n426_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G113gat), .B(G120gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n429_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n439_), .B(KEYINPUT31), .Z(new_n440_));
  NAND3_X1  g239(.A1(new_n417_), .A2(new_n423_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n421_), .A2(KEYINPUT84), .A3(new_n422_), .A4(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G1gat), .B(G29gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(new_n242_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT0), .B(G57gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT3), .ZN(new_n449_));
  INV_X1    g248(.A(G141gat), .ZN(new_n450_));
  INV_X1    g249(.A(G148gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G141gat), .A2(G148gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT2), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n452_), .A2(new_n455_), .A3(new_n456_), .A4(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT85), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(G155gat), .A2(G162gat), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT85), .B1(new_n464_), .B2(new_n459_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n458_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n459_), .A2(KEYINPUT1), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT1), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G155gat), .A3(G162gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n469_), .A3(new_n464_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n450_), .A2(new_n451_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n453_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n466_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n438_), .A3(new_n437_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n429_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n435_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n466_), .B(new_n472_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n477_), .A3(KEYINPUT4), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT4), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n473_), .A2(new_n479_), .A3(new_n438_), .A4(new_n437_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G225gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT94), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n474_), .A2(new_n477_), .A3(new_n481_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n448_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n485_), .A3(new_n448_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G228gat), .A2(G233gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G197gat), .B(G204gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT21), .ZN(new_n495_));
  INV_X1    g294(.A(G211gat), .ZN(new_n496_));
  INV_X1    g295(.A(G218gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G211gat), .A2(G218gat), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n494_), .A2(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT90), .B1(new_n494_), .B2(new_n495_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502_));
  INV_X1    g301(.A(G204gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G197gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n503_), .A2(G197gat), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n502_), .B(KEYINPUT21), .C1(new_n505_), .C2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n500_), .A2(new_n501_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G197gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(G204gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n504_), .A2(new_n510_), .A3(new_n495_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n498_), .A2(new_n499_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT21), .B1(new_n505_), .B2(new_n506_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT90), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n508_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n493_), .B1(new_n516_), .B2(KEYINPUT88), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G78gat), .B(G106gat), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n508_), .A2(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n473_), .A2(KEYINPUT29), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT29), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n466_), .B2(new_n472_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n518_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n516_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n517_), .B1(new_n521_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n519_), .A2(new_n520_), .A3(new_n518_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n516_), .B2(new_n523_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT88), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n519_), .A2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n528_), .A2(new_n529_), .A3(new_n531_), .A4(new_n493_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n526_), .A2(new_n527_), .A3(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n466_), .A2(new_n522_), .A3(new_n472_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G22gat), .B(G50gat), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n534_), .B(new_n535_), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n538_));
  INV_X1    g337(.A(new_n536_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n526_), .A2(new_n539_), .A3(new_n527_), .A4(new_n532_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n537_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT27), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n392_), .A2(new_n403_), .A3(new_n516_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n402_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n382_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT92), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n396_), .A2(new_n548_), .A3(new_n383_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n396_), .B2(new_n383_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n388_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n389_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT91), .B1(new_n390_), .B2(new_n388_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n400_), .A2(new_n399_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n374_), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT80), .B1(G183gat), .B2(G190gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT23), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n556_), .A2(new_n387_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n547_), .A2(new_n551_), .B1(new_n561_), .B2(new_n386_), .ZN(new_n562_));
  OAI211_X1 g361(.A(KEYINPUT20), .B(new_n545_), .C1(new_n562_), .C2(new_n516_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G226gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT19), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G64gat), .B(G92gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(G8gat), .B(G36gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n392_), .A2(new_n403_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n519_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n565_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n562_), .A2(new_n516_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n566_), .A2(new_n572_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n572_), .B1(new_n566_), .B2(new_n578_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n544_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n563_), .A2(new_n565_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n576_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n571_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n566_), .A2(new_n572_), .A3(new_n578_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(KEYINPUT27), .A3(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n444_), .A2(new_n490_), .A3(new_n543_), .A4(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n579_), .A2(new_n580_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n478_), .A2(new_n481_), .A3(new_n480_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n448_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n474_), .A2(new_n477_), .A3(new_n483_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT95), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n488_), .B(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n589_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n572_), .A2(KEYINPUT32), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n566_), .A2(new_n578_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n488_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n600_), .B1(new_n601_), .B2(new_n486_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n563_), .A2(new_n565_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n583_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n599_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n598_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(KEYINPUT32), .B(new_n572_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n489_), .A2(new_n607_), .A3(KEYINPUT96), .A4(new_n600_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n597_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n541_), .A2(new_n542_), .A3(new_n489_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n609_), .A2(new_n543_), .B1(new_n610_), .B2(new_n587_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n588_), .B1(new_n611_), .B2(new_n444_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n367_), .B(new_n612_), .C1(KEYINPUT76), .C2(new_n366_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT97), .Z(new_n614_));
  XOR2_X1   g413(.A(new_n489_), .B(KEYINPUT98), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(new_n203_), .A3(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n313_), .A2(new_n228_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n609_), .A2(new_n543_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n610_), .A2(new_n587_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n444_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n620_), .B1(new_n625_), .B2(new_n588_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n349_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n365_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G1gat), .B1(new_n629_), .B2(new_n490_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n619_), .A2(new_n630_), .ZN(G1324gat));
  INV_X1    g430(.A(new_n587_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n614_), .A2(new_n204_), .A3(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G8gat), .B1(new_n629_), .B2(new_n587_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT39), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1325gat));
  OAI21_X1  g437(.A(G15gat), .B1(new_n629_), .B2(new_n624_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT41), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n613_), .A2(G15gat), .A3(new_n624_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1326gat));
  OAI21_X1  g441(.A(G22gat), .B1(new_n629_), .B2(new_n543_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT42), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n613_), .A2(G22gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(new_n543_), .ZN(G1327gat));
  INV_X1    g445(.A(new_n365_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n349_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n626_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n489_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n349_), .B(KEYINPUT37), .C1(KEYINPUT72), .C2(new_n338_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n338_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n339_), .A2(new_n654_), .A3(new_n344_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n625_), .B2(new_n588_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n651_), .B(new_n652_), .C1(new_n657_), .C2(KEYINPUT101), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT101), .B1(new_n612_), .B2(new_n350_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT43), .B1(new_n659_), .B2(KEYINPUT102), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n612_), .A2(new_n350_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT102), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(new_n660_), .A3(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n647_), .A2(new_n620_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT104), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(new_n664_), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT104), .B1(new_n665_), .B2(KEYINPUT103), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n668_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n663_), .A2(new_n664_), .A3(new_n666_), .A4(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(new_n615_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n650_), .B1(new_n674_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n649_), .A2(new_n676_), .A3(new_n632_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT45), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n672_), .B2(new_n632_), .ZN(new_n681_));
  AOI211_X1 g480(.A(KEYINPUT105), .B(new_n587_), .C1(new_n669_), .C2(new_n671_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n679_), .B1(new_n683_), .B2(G36gat), .ZN(new_n684_));
  NOR4_X1   g483(.A1(new_n681_), .A2(new_n682_), .A3(KEYINPUT106), .A4(new_n676_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n678_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT107), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n687_), .A2(KEYINPUT107), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n686_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n672_), .A2(new_n632_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT105), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n672_), .A2(new_n680_), .A3(new_n632_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(G36gat), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT106), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n683_), .A2(new_n679_), .A3(G36gat), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n697_), .A2(KEYINPUT107), .A3(new_n687_), .A4(new_n678_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n690_), .A2(new_n698_), .ZN(G1329gat));
  NAND3_X1  g498(.A1(new_n672_), .A2(G43gat), .A3(new_n444_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT108), .Z(new_n701_));
  AND2_X1   g500(.A1(new_n649_), .A2(new_n444_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT109), .B(G43gat), .Z(new_n703_));
  OAI21_X1  g502(.A(new_n701_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g504(.A(G50gat), .B1(new_n673_), .B2(new_n543_), .ZN(new_n706_));
  INV_X1    g505(.A(G50gat), .ZN(new_n707_));
  INV_X1    g506(.A(new_n543_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n649_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(G1331gat));
  NOR2_X1   g509(.A1(new_n313_), .A2(new_n228_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n612_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n628_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n713_), .A2(new_n270_), .A3(new_n490_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n712_), .A2(new_n647_), .A3(new_n656_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n616_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n716_), .B2(new_n270_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n713_), .B2(new_n587_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT48), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n715_), .A2(new_n271_), .A3(new_n632_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n713_), .B2(new_n624_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n715_), .A2(new_n407_), .A3(new_n444_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1334gat));
  OAI21_X1  g524(.A(G78gat), .B1(new_n713_), .B2(new_n543_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT50), .ZN(new_n727_));
  INV_X1    g526(.A(G78gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n715_), .A2(new_n728_), .A3(new_n708_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT110), .Z(G1335gat));
  NAND3_X1  g530(.A1(new_n663_), .A2(new_n365_), .A3(new_n711_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT111), .Z(new_n733_));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n490_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n712_), .A2(new_n648_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n242_), .A3(new_n616_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1336gat));
  OAI21_X1  g536(.A(G92gat), .B1(new_n733_), .B2(new_n587_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n735_), .A2(new_n243_), .A3(new_n632_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1337gat));
  OAI21_X1  g539(.A(G99gat), .B1(new_n732_), .B2(new_n624_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n624_), .A2(new_n257_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n735_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g544(.A(G106gat), .B1(new_n732_), .B2(new_n543_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n747_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(KEYINPUT52), .A3(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n735_), .A2(new_n232_), .A3(new_n708_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n747_), .A3(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n751_), .A3(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(G1339gat));
  AOI21_X1  g555(.A(new_n295_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n298_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n294_), .A2(new_n297_), .A3(KEYINPUT55), .A4(new_n295_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n305_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT56), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(new_n764_), .A3(new_n305_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n763_), .A2(new_n228_), .A3(new_n307_), .A4(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT114), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n764_), .B1(new_n761_), .B2(new_n305_), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT56), .B(new_n304_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n228_), .A4(new_n307_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n219_), .A2(new_n217_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n227_), .B1(new_n216_), .B2(new_n220_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n223_), .A2(new_n227_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n308_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n767_), .A2(new_n772_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT57), .B1(new_n777_), .B2(new_n349_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n763_), .A2(new_n307_), .A3(new_n775_), .A4(new_n765_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT58), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n770_), .A2(KEYINPUT58), .A3(new_n307_), .A4(new_n775_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n350_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n778_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n777_), .A2(KEYINPUT57), .A3(new_n349_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n647_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n366_), .A2(new_n229_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT54), .Z(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n444_), .A2(new_n616_), .A3(new_n543_), .A4(new_n587_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(G113gat), .B1(new_n792_), .B2(new_n228_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT115), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n795_));
  XOR2_X1   g594(.A(new_n791_), .B(KEYINPUT117), .Z(new_n796_));
  INV_X1    g595(.A(new_n786_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n785_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT118), .B1(new_n778_), .B2(new_n784_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n647_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n795_), .B(new_n796_), .C1(new_n801_), .C2(new_n789_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT119), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n777_), .A2(new_n349_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n798_), .A3(new_n783_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(new_n786_), .A3(new_n800_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n789_), .B1(new_n808_), .B2(new_n365_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n810_), .A2(new_n811_), .A3(new_n795_), .A4(new_n796_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n803_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT59), .B1(new_n790_), .B2(new_n791_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n228_), .A2(G113gat), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT120), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n794_), .B1(new_n815_), .B2(new_n817_), .ZN(G1340gat));
  INV_X1    g617(.A(G120gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n313_), .B2(KEYINPUT60), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n792_), .B(new_n820_), .C1(KEYINPUT60), .C2(new_n819_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n815_), .A2(new_n314_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n819_), .ZN(G1341gat));
  AOI21_X1  g622(.A(G127gat), .B1(new_n792_), .B2(new_n647_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n815_), .A2(G127gat), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n647_), .ZN(G1342gat));
  NAND4_X1  g625(.A1(new_n813_), .A2(new_n814_), .A3(G134gat), .A4(new_n350_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n790_), .A2(new_n349_), .A3(new_n791_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n828_), .A2(G134gat), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n827_), .A2(KEYINPUT121), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1343gat));
  NOR3_X1   g633(.A1(new_n790_), .A2(new_n543_), .A3(new_n444_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n632_), .A2(new_n615_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n229_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(new_n450_), .ZN(G1344gat));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n313_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(new_n451_), .ZN(G1345gat));
  NOR2_X1   g640(.A1(new_n837_), .A2(new_n365_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT61), .B(G155gat), .Z(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1346gat));
  INV_X1    g643(.A(new_n837_), .ZN(new_n845_));
  AOI21_X1  g644(.A(G162gat), .B1(new_n845_), .B2(new_n627_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n350_), .A2(G162gat), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT122), .Z(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n845_), .B2(new_n848_), .ZN(G1347gat));
  NOR3_X1   g648(.A1(new_n624_), .A2(new_n616_), .A3(new_n587_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n809_), .A2(new_n229_), .A3(new_n708_), .A4(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(G169gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT123), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n543_), .B(new_n850_), .C1(new_n801_), .C2(new_n789_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n855_), .B(G169gat), .C1(new_n856_), .C2(new_n229_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(KEYINPUT62), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n852_), .B1(new_n395_), .B2(new_n394_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT123), .B(new_n860_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n858_), .A2(new_n859_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT124), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n858_), .A2(new_n864_), .A3(new_n859_), .A4(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1348gat));
  OAI21_X1  g665(.A(new_n393_), .B1(new_n856_), .B2(new_n313_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n790_), .A2(new_n708_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n868_), .A2(G176gat), .A3(new_n850_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n313_), .B2(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT125), .ZN(G1349gat));
  NOR2_X1   g670(.A1(new_n851_), .A2(new_n365_), .ZN(new_n872_));
  AOI21_X1  g671(.A(G183gat), .B1(new_n868_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n856_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n365_), .A2(new_n556_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT126), .ZN(G1350gat));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n627_), .A3(new_n387_), .ZN(new_n878_));
  OAI21_X1  g677(.A(G190gat), .B1(new_n856_), .B2(new_n656_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1351gat));
  NOR2_X1   g679(.A1(new_n790_), .A2(new_n444_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n610_), .A3(new_n632_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n229_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n509_), .ZN(G1352gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n313_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n503_), .ZN(G1353gat));
  NOR2_X1   g685(.A1(new_n882_), .A2(new_n365_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT63), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n496_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n887_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT127), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT127), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n887_), .A2(new_n893_), .A3(new_n890_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n888_), .A2(new_n496_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n892_), .A2(new_n888_), .A3(new_n496_), .A4(new_n894_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1354gat));
  NOR3_X1   g698(.A1(new_n882_), .A2(new_n497_), .A3(new_n656_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n882_), .A2(new_n349_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n497_), .B2(new_n901_), .ZN(G1355gat));
endmodule


