//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_;
  INV_X1    g000(.A(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT26), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT77), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  AND2_X1   g004(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G190gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n203_), .A2(new_n210_), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n205_), .B(new_n208_), .C1(new_n211_), .C2(new_n204_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(new_n202_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n212_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n215_), .B(new_n216_), .C1(G183gat), .C2(G190gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n227_), .A3(new_n221_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT78), .ZN(new_n230_));
  XOR2_X1   g029(.A(G71gat), .B(G99gat), .Z(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT30), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n230_), .B(new_n232_), .Z(new_n233_));
  XNOR2_X1  g032(.A(G15gat), .B(G43gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n235_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239_));
  INV_X1    g038(.A(G113gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G120gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT80), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(KEYINPUT80), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT31), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT31), .B1(new_n244_), .B2(new_n245_), .ZN(new_n249_));
  OR3_X1    g048(.A1(new_n248_), .A2(KEYINPUT79), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G227gat), .A2(G233gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n250_), .A2(new_n252_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n238_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n250_), .A2(new_n252_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n257_), .A2(new_n253_), .A3(new_n236_), .A4(new_n237_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G78gat), .B(G106gat), .Z(new_n260_));
  INV_X1    g059(.A(G204gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(G197gat), .ZN(new_n262_));
  INV_X1    g061(.A(G197gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT87), .B1(new_n263_), .B2(G204gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(new_n261_), .A3(G197gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n262_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268_));
  OR2_X1    g067(.A1(G211gat), .A2(G218gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G211gat), .A2(G218gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n267_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n263_), .A2(G204gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n261_), .A2(G197gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n276_), .A2(KEYINPUT21), .B1(new_n269_), .B2(new_n270_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n265_), .B1(G197gat), .B2(new_n261_), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n263_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n268_), .B(new_n274_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT88), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n277_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n273_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT81), .ZN(new_n285_));
  INV_X1    g084(.A(G155gat), .ZN(new_n286_));
  INV_X1    g085(.A(G162gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT84), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n294_));
  NOR2_X1   g093(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT3), .ZN(new_n299_));
  INV_X1    g098(.A(G141gat), .ZN(new_n300_));
  INV_X1    g099(.A(G148gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(KEYINPUT83), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n297_), .A2(new_n298_), .A3(new_n302_), .A4(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n288_), .A2(KEYINPUT84), .A3(new_n289_), .A4(new_n290_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n293_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n293_), .A2(new_n304_), .A3(KEYINPUT85), .A4(new_n305_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n290_), .A2(KEYINPUT1), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(G155gat), .A3(G162gat), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n288_), .A2(new_n310_), .A3(new_n312_), .A4(new_n289_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n300_), .A2(new_n301_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n314_), .A3(new_n296_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n313_), .A2(KEYINPUT82), .A3(new_n314_), .A4(new_n296_), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n308_), .A2(new_n309_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n284_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(G228gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(G228gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n323_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n322_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n330_), .B(new_n284_), .C1(new_n319_), .C2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n260_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT90), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n319_), .A2(new_n331_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G22gat), .B(G50gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT28), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n336_), .B(new_n339_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n329_), .A2(new_n260_), .A3(new_n332_), .ZN(new_n341_));
  OAI22_X1  g140(.A1(new_n335_), .A2(new_n340_), .B1(new_n341_), .B2(new_n333_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n308_), .A2(new_n309_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n317_), .A2(new_n318_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n328_), .B1(new_n345_), .B2(KEYINPUT29), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n346_), .A2(new_n284_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n260_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n329_), .A2(new_n332_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n260_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n340_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n348_), .A2(new_n351_), .A3(new_n352_), .A4(new_n334_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n342_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT18), .B(G64gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G92gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n203_), .B(new_n210_), .C1(new_n206_), .C2(new_n207_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n222_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT91), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(KEYINPUT91), .A3(new_n222_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n220_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n228_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT92), .B1(new_n284_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n228_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n360_), .A2(KEYINPUT91), .A3(new_n222_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT91), .B1(new_n360_), .B2(new_n222_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n371_), .B2(new_n220_), .ZN(new_n372_));
  AOI211_X1 g171(.A(KEYINPUT21), .B(new_n262_), .C1(new_n264_), .C2(new_n266_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G197gat), .B(G204gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n271_), .B1(new_n374_), .B2(new_n268_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT88), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n277_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n272_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT92), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n372_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n367_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n284_), .A2(new_n229_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G226gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT19), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(KEYINPUT20), .A3(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n381_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n284_), .B2(new_n366_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n378_), .A2(new_n228_), .A3(new_n223_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n385_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n359_), .B1(new_n387_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n393_));
  INV_X1    g192(.A(new_n391_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n384_), .B1(new_n284_), .B2(new_n229_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n367_), .A2(new_n395_), .A3(new_n380_), .A4(KEYINPUT20), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n396_), .A3(new_n358_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n392_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n387_), .A2(new_n391_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(KEYINPUT93), .A3(new_n358_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G1gat), .B(G29gat), .Z(new_n402_));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n404_), .B(new_n405_), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT94), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n343_), .A2(new_n408_), .A3(new_n344_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n243_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n319_), .A2(new_n408_), .A3(new_n243_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(KEYINPUT4), .A3(new_n414_), .ZN(new_n416_));
  OR3_X1    g215(.A1(new_n319_), .A2(KEYINPUT4), .A3(new_n243_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n407_), .B(new_n415_), .C1(new_n418_), .C2(new_n413_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT33), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n413_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n413_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n420_), .B1(new_n424_), .B2(new_n406_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n412_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n420_), .B(new_n406_), .C1(new_n426_), .C2(new_n422_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n401_), .B(new_n419_), .C1(new_n425_), .C2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n358_), .A2(KEYINPUT32), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n382_), .B(KEYINPUT20), .C1(new_n284_), .C2(new_n366_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n384_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n389_), .A2(new_n390_), .A3(new_n385_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n430_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT97), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n430_), .B(KEYINPUT96), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n399_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n421_), .A2(new_n407_), .A3(new_n423_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n406_), .B1(new_n426_), .B2(new_n422_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n435_), .B(new_n437_), .C1(new_n439_), .C2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n354_), .B1(new_n429_), .B2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n438_), .A2(new_n440_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT27), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n398_), .A2(new_n446_), .A3(new_n400_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n432_), .A2(new_n433_), .ZN(new_n448_));
  OAI211_X1 g247(.A(KEYINPUT27), .B(new_n397_), .C1(new_n448_), .C2(new_n358_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT90), .B1(new_n347_), .B2(new_n260_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n451_), .A2(new_n352_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n452_));
  NOR4_X1   g251(.A1(new_n341_), .A2(new_n333_), .A3(new_n340_), .A4(KEYINPUT90), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n445_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n259_), .B1(new_n443_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT98), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT98), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n458_), .B(new_n259_), .C1(new_n443_), .C2(new_n455_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT99), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n450_), .B2(new_n354_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n454_), .A2(KEYINPUT99), .A3(new_n447_), .A4(new_n449_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n445_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT100), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT100), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n457_), .A2(new_n459_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT13), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G230gat), .A2(G233gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G99gat), .A2(G106gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT6), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT10), .B(G99gat), .ZN(new_n475_));
  INV_X1    g274(.A(G85gat), .ZN(new_n476_));
  INV_X1    g275(.A(G92gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT64), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT9), .ZN(new_n479_));
  NOR2_X1   g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  OAI221_X1 g279(.A(new_n474_), .B1(G106gat), .B2(new_n475_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT8), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT7), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n483_), .B1(KEYINPUT65), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT65), .B(KEYINPUT7), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n483_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT66), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT66), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n489_), .B(new_n485_), .C1(new_n486_), .C2(new_n483_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n474_), .A3(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G85gat), .B(G92gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n482_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n487_), .ZN(new_n495_));
  AOI211_X1 g294(.A(KEYINPUT8), .B(new_n492_), .C1(new_n495_), .C2(new_n474_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n481_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G71gat), .B(G78gat), .ZN(new_n501_));
  OR3_X1    g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n501_), .A3(KEYINPUT11), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n497_), .A2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n506_), .A2(KEYINPUT12), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n481_), .B(new_n504_), .C1(new_n494_), .C2(new_n496_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(KEYINPUT12), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n472_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n471_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT67), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n511_), .A2(KEYINPUT67), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G120gat), .B(G148gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(new_n261_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT5), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(new_n226_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n512_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n470_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(KEYINPUT13), .A3(new_n522_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(G141gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT74), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n240_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531_));
  INV_X1    g330(.A(G1gat), .ZN(new_n532_));
  INV_X1    g331(.A(G8gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT14), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G1gat), .B(G8gat), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n536_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT15), .ZN(new_n541_));
  XOR2_X1   g340(.A(G29gat), .B(G36gat), .Z(new_n542_));
  INV_X1    g341(.A(G43gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G29gat), .B(G36gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(G43gat), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n544_), .A2(G50gat), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(G50gat), .B1(new_n544_), .B2(new_n546_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n547_), .A2(new_n548_), .A3(KEYINPUT69), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT69), .ZN(new_n550_));
  INV_X1    g349(.A(G50gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n546_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n545_), .A2(G43gat), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n544_), .A2(G50gat), .A3(new_n546_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n550_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n541_), .B1(new_n549_), .B2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT69), .B1(new_n547_), .B2(new_n548_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(new_n550_), .A3(new_n555_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(KEYINPUT15), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n540_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n554_), .A2(new_n538_), .A3(new_n537_), .A4(new_n555_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n562_), .A2(KEYINPUT72), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(KEYINPUT72), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n561_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT73), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n547_), .A2(new_n548_), .ZN(new_n570_));
  OAI22_X1  g369(.A1(new_n563_), .A2(new_n564_), .B1(new_n540_), .B2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n571_), .B2(new_n567_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n557_), .A2(new_n560_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n539_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n563_), .A2(new_n564_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n575_), .A2(KEYINPUT73), .A3(new_n566_), .A4(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n530_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n577_), .B(new_n530_), .C1(new_n568_), .C2(new_n572_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT76), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n580_), .A2(KEYINPUT75), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n580_), .B2(KEYINPUT75), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n579_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(KEYINPUT75), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT76), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n580_), .A2(KEYINPUT75), .A3(new_n581_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n578_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n469_), .A2(new_n526_), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(G134gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(new_n287_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT35), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT68), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT34), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n574_), .A2(new_n497_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n481_), .B(new_n570_), .C1(new_n494_), .C2(new_n496_), .ZN(new_n604_));
  AOI211_X1 g403(.A(new_n598_), .B(new_n602_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(KEYINPUT35), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n598_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .A4(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n596_), .B(new_n597_), .C1(new_n605_), .C2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n603_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(KEYINPUT35), .A3(new_n601_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n595_), .A3(new_n608_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n610_), .A2(new_n613_), .A3(KEYINPUT70), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n504_), .B(new_n540_), .ZN(new_n617_));
  AND2_X1   g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT16), .B(G183gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(G211gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(KEYINPUT71), .A3(KEYINPUT17), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(KEYINPUT17), .B2(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n619_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n610_), .A2(new_n613_), .A3(KEYINPUT70), .A4(KEYINPUT37), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n616_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n590_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n532_), .A3(new_n445_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT38), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n610_), .A2(new_n613_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n629_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n590_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n639_), .B2(new_n444_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n634_), .A2(new_n640_), .ZN(G1324gat));
  INV_X1    g440(.A(new_n450_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G8gat), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(KEYINPUT101), .B(G8gat), .C1(new_n639_), .C2(new_n642_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(KEYINPUT39), .A3(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n632_), .A2(new_n533_), .A3(new_n450_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n643_), .A2(new_n644_), .A3(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n639_), .B2(new_n259_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT41), .Z(new_n655_));
  INV_X1    g454(.A(G15gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n259_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n632_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(G1326gat));
  OAI21_X1  g458(.A(G22gat), .B1(new_n639_), .B2(new_n454_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n632_), .A2(new_n662_), .A3(new_n354_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1327gat));
  NAND2_X1  g463(.A1(new_n457_), .A2(new_n459_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n466_), .A2(new_n468_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n636_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n526_), .A2(new_n589_), .A3(new_n629_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G29gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n445_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n616_), .A2(new_n630_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n469_), .B2(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n469_), .A2(KEYINPUT43), .A3(new_n677_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT103), .B(new_n675_), .C1(new_n469_), .C2(new_n677_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT44), .B(new_n670_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n677_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n680_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n687_), .A2(new_n674_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n682_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n686_), .B1(new_n691_), .B2(new_n669_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n444_), .B1(new_n684_), .B2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n673_), .B1(new_n694_), .B2(new_n672_), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n696_), .A2(KEYINPUT105), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT106), .Z(new_n698_));
  OAI21_X1  g497(.A(new_n450_), .B1(new_n683_), .B2(new_n692_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n701_));
  INV_X1    g500(.A(G36gat), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n671_), .A2(new_n701_), .A3(new_n702_), .A4(new_n450_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n469_), .A2(new_n635_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(new_n702_), .A3(new_n669_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT45), .B1(new_n705_), .B2(new_n642_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n696_), .A2(KEYINPUT105), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n698_), .B1(new_n700_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n698_), .ZN(new_n712_));
  AOI211_X1 g511(.A(new_n712_), .B(new_n709_), .C1(new_n699_), .C2(G36gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1329gat));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n657_), .B1(new_n683_), .B2(new_n692_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G43gat), .ZN(new_n717_));
  NOR4_X1   g516(.A1(new_n668_), .A2(G43gat), .A3(new_n259_), .A4(new_n670_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n715_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT47), .B(new_n718_), .C1(new_n716_), .C2(G43gat), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1330gat));
  NAND3_X1  g521(.A1(new_n671_), .A2(new_n551_), .A3(new_n354_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n454_), .B1(new_n684_), .B2(new_n693_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n551_), .ZN(G1331gat));
  INV_X1    g524(.A(new_n526_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n584_), .A2(new_n588_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n469_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n728_), .A2(G57gat), .A3(new_n445_), .A4(new_n638_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT107), .Z(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n631_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n445_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1332gat));
  NAND2_X1  g533(.A1(new_n728_), .A2(new_n638_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G64gat), .B1(new_n735_), .B2(new_n642_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT48), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n642_), .A2(G64gat), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT108), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n737_), .B1(new_n731_), .B2(new_n739_), .ZN(G1333gat));
  OAI21_X1  g539(.A(G71gat), .B1(new_n735_), .B2(new_n259_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT49), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n259_), .A2(G71gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n731_), .B2(new_n743_), .ZN(G1334gat));
  OAI21_X1  g543(.A(G78gat), .B1(new_n735_), .B2(new_n454_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT50), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n454_), .A2(G78gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n731_), .B2(new_n747_), .ZN(G1335gat));
  NOR3_X1   g547(.A1(new_n726_), .A2(new_n727_), .A3(new_n629_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n704_), .A2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT109), .Z(new_n751_));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n445_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n691_), .A2(new_n749_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(new_n445_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(G85gat), .B2(new_n754_), .ZN(G1336gat));
  AOI21_X1  g554(.A(G92gat), .B1(new_n751_), .B2(new_n450_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n642_), .A2(new_n477_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n753_), .B2(new_n757_), .ZN(G1337gat));
  INV_X1    g557(.A(new_n475_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n751_), .A2(new_n759_), .A3(new_n657_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n691_), .A2(new_n657_), .A3(new_n749_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(G99gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(G99gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT51), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n760_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1338gat));
  INV_X1    g568(.A(G106gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n751_), .A2(new_n770_), .A3(new_n354_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n691_), .A2(new_n354_), .A3(new_n749_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(new_n773_), .A3(G106gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n772_), .B2(G106gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n771_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n657_), .A2(new_n445_), .A3(new_n463_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n510_), .B(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n507_), .A2(new_n472_), .A3(new_n509_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n518_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n522_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n575_), .A2(new_n567_), .A3(new_n576_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n530_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n571_), .A2(new_n566_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n794_), .A2(KEYINPUT113), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(KEYINPUT113), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n580_), .A3(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n507_), .A2(new_n509_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n785_), .B1(new_n798_), .B2(new_n472_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n510_), .A2(KEYINPUT55), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n787_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n519_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n797_), .B1(new_n802_), .B2(KEYINPUT56), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n784_), .B1(new_n790_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n523_), .B1(new_n802_), .B2(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n788_), .A2(new_n789_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT58), .A4(new_n797_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n804_), .A2(new_n676_), .A3(new_n807_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n809_));
  OAI21_X1  g608(.A(new_n797_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT112), .B1(new_n789_), .B2(KEYINPUT111), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n789_), .A2(KEYINPUT112), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n801_), .A2(new_n519_), .A3(new_n812_), .A4(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(new_n584_), .A3(new_n522_), .A4(new_n588_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n802_), .A2(new_n811_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n810_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n809_), .B1(new_n818_), .B2(new_n635_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n808_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(KEYINPUT57), .A3(new_n635_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n629_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n631_), .A2(new_n524_), .A3(new_n525_), .A4(new_n589_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n783_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n781_), .B1(new_n826_), .B2(KEYINPUT59), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n804_), .A2(new_n676_), .A3(new_n807_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n727_), .A2(new_n522_), .A3(new_n816_), .A4(new_n814_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n636_), .B1(new_n829_), .B2(new_n810_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n821_), .B(new_n828_), .C1(new_n830_), .C2(new_n809_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n825_), .B1(new_n831_), .B2(new_n637_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n781_), .B(KEYINPUT59), .C1(new_n832_), .C2(new_n782_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n827_), .A2(new_n834_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n836_));
  INV_X1    g635(.A(new_n821_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n828_), .B1(new_n830_), .B2(new_n809_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(KEYINPUT117), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n820_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n629_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n783_), .B(new_n836_), .C1(new_n842_), .C2(new_n825_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n835_), .A2(G113gat), .A3(new_n727_), .A4(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n240_), .B1(new_n826_), .B2(new_n589_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1340gat));
  NAND4_X1  g645(.A1(new_n835_), .A2(KEYINPUT118), .A3(new_n526_), .A4(new_n843_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n843_), .B(new_n526_), .C1(new_n827_), .C2(new_n834_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(G120gat), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n826_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n242_), .B1(new_n726_), .B2(KEYINPUT60), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n852_), .B(new_n853_), .C1(KEYINPUT60), .C2(new_n242_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(G1341gat));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n843_), .B(new_n629_), .C1(new_n827_), .C2(new_n834_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G127gat), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n826_), .A2(G127gat), .A3(new_n637_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n856_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  AOI211_X1 g660(.A(KEYINPUT119), .B(new_n859_), .C1(new_n857_), .C2(G127gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1342gat));
  AOI21_X1  g662(.A(G134gat), .B1(new_n852_), .B2(new_n636_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n835_), .A2(new_n676_), .A3(new_n843_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g665(.A1(new_n259_), .A2(new_n354_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n832_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n450_), .A2(new_n444_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT120), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n868_), .A2(new_n872_), .A3(new_n869_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n727_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n526_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT121), .B(G148gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1345gat));
  NAND2_X1  g678(.A1(new_n874_), .A2(new_n629_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT61), .B(G155gat), .Z(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT122), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n880_), .B(new_n882_), .ZN(G1346gat));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n635_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(G162gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n676_), .A2(G162gat), .ZN(new_n887_));
  XOR2_X1   g686(.A(new_n887_), .B(KEYINPUT123), .Z(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n884_), .B1(new_n886_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n890_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n892_), .B(KEYINPUT124), .C1(G162gat), .C2(new_n885_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1347gat));
  OR2_X1    g693(.A1(new_n842_), .A2(new_n825_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n464_), .A2(new_n450_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n895_), .A2(new_n727_), .A3(new_n454_), .A4(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n897_), .A2(new_n898_), .A3(G169gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n897_), .B2(G169gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n895_), .A2(new_n454_), .A3(new_n896_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n727_), .A2(new_n225_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT125), .ZN(new_n903_));
  OAI22_X1  g702(.A1(new_n899_), .A2(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(G1348gat));
  INV_X1    g703(.A(new_n901_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G176gat), .B1(new_n905_), .B2(new_n526_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n832_), .A2(new_n354_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n896_), .A2(new_n526_), .A3(G176gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1349gat));
  NOR3_X1   g708(.A1(new_n901_), .A2(new_n208_), .A3(new_n637_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n896_), .A2(new_n629_), .ZN(new_n911_));
  AOI21_X1  g710(.A(G183gat), .B1(new_n907_), .B2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n901_), .B2(new_n677_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n636_), .A2(new_n211_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n901_), .B2(new_n915_), .ZN(G1351gat));
  NOR2_X1   g715(.A1(new_n642_), .A2(new_n445_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n868_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n589_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT127), .B1(new_n919_), .B2(KEYINPUT126), .ZN(new_n920_));
  AOI21_X1  g719(.A(G197gat), .B1(new_n919_), .B2(KEYINPUT126), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n922_), .B(new_n923_), .C1(new_n918_), .C2(new_n589_), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n920_), .A2(new_n921_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n921_), .B1(new_n924_), .B2(new_n920_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1352gat));
  NOR2_X1   g726(.A1(new_n918_), .A2(new_n726_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(new_n261_), .ZN(G1353gat));
  INV_X1    g728(.A(new_n918_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n629_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  AND2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n931_), .B2(new_n932_), .ZN(G1354gat));
  NOR2_X1   g734(.A1(new_n918_), .A2(new_n635_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n930_), .A2(new_n676_), .ZN(new_n937_));
  MUX2_X1   g736(.A(new_n936_), .B(new_n937_), .S(G218gat), .Z(G1355gat));
endmodule


