//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT36), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G232gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT34), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT35), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT68), .Z(new_n210_));
  INV_X1    g009(.A(KEYINPUT72), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n212_), .B(KEYINPUT6), .Z(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n213_), .B1(new_n218_), .B2(KEYINPUT66), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(KEYINPUT66), .B2(new_n218_), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  INV_X1    g020(.A(G92gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n220_), .A2(KEYINPUT8), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G29gat), .B(G36gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n227_), .A2(KEYINPUT69), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(KEYINPUT69), .ZN(new_n229_));
  XOR2_X1   g028(.A(G43gat), .B(G50gat), .Z(new_n230_));
  OR3_X1    g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n224_), .B1(new_n223_), .B2(KEYINPUT9), .ZN(new_n234_));
  INV_X1    g033(.A(new_n223_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT9), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n235_), .A2(KEYINPUT64), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT64), .B1(new_n235_), .B2(new_n236_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n234_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G106gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT10), .B(G99gat), .Z(new_n241_));
  AOI21_X1  g040(.A(new_n213_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n225_), .B1(new_n218_), .B2(new_n213_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT8), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n239_), .A2(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n226_), .A2(new_n233_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n226_), .A2(KEYINPUT71), .A3(new_n233_), .A4(new_n245_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n208_), .A2(KEYINPUT35), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n211_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n226_), .A2(new_n245_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT15), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT15), .B1(new_n231_), .B2(new_n232_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n253_), .A2(new_n256_), .A3(KEYINPUT70), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT70), .B1(new_n253_), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n259_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n248_), .A2(new_n251_), .A3(new_n211_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n210_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n248_), .A2(new_n251_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n210_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n206_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n204_), .A2(new_n205_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n262_), .A2(new_n265_), .A3(new_n205_), .A4(new_n204_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT37), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n268_), .A2(new_n269_), .A3(KEYINPUT37), .A4(new_n270_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G57gat), .B(G64gat), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(KEYINPUT11), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(KEYINPUT11), .ZN(new_n278_));
  XOR2_X1   g077(.A(G71gat), .B(G78gat), .Z(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n278_), .A2(new_n279_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n253_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n226_), .A2(new_n282_), .A3(new_n245_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G230gat), .ZN(new_n287_));
  INV_X1    g086(.A(G233gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT67), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT67), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(new_n292_), .A3(new_n289_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n284_), .A2(KEYINPUT12), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n284_), .A2(KEYINPUT12), .A3(new_n285_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n289_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G120gat), .B(G148gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT5), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G176gat), .B(G204gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n294_), .A2(new_n298_), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n294_), .B2(new_n298_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT13), .ZN(new_n306_));
  OR3_X1    g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n306_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G231gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n282_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT74), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G15gat), .B(G22gat), .ZN(new_n314_));
  INV_X1    g113(.A(G1gat), .ZN(new_n315_));
  INV_X1    g114(.A(G8gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT14), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G1gat), .B(G8gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n313_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G127gat), .B(G155gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT16), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G183gat), .B(G211gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT17), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n327_), .A2(new_n328_), .ZN(new_n330_));
  OR3_X1    g129(.A1(new_n323_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n323_), .A2(new_n329_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n275_), .A2(new_n310_), .A3(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G8gat), .B(G36gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT93), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT88), .ZN(new_n344_));
  XOR2_X1   g143(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(G204gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT85), .B1(new_n347_), .B2(G197gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349_));
  INV_X1    g148(.A(G197gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(G204gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(G197gat), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n348_), .A2(new_n351_), .A3(KEYINPUT86), .A4(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT21), .ZN(new_n354_));
  INV_X1    g153(.A(G218gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G211gat), .ZN(new_n356_));
  INV_X1    g155(.A(G211gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G218gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n354_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n348_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT86), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n348_), .A2(new_n351_), .A3(new_n354_), .A4(new_n352_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n356_), .A2(new_n358_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n350_), .A2(G204gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n352_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(KEYINPUT21), .B2(new_n367_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n360_), .A2(new_n363_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G190gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT26), .B1(new_n370_), .B2(KEYINPUT77), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT26), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(G190gat), .ZN(new_n374_));
  INV_X1    g173(.A(G183gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT25), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G183gat), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n371_), .A2(new_n374_), .A3(new_n376_), .A4(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT25), .B(G183gat), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n382_), .A2(KEYINPUT78), .A3(new_n371_), .A4(new_n374_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G169gat), .ZN(new_n385_));
  INV_X1    g184(.A(G176gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(KEYINPUT24), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT23), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(G183gat), .A3(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  OR3_X1    g193(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n389_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n384_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT80), .B1(new_n385_), .B2(KEYINPUT22), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT22), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(G169gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n401_), .A3(new_n386_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT22), .B1(KEYINPUT79), .B2(G169gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(KEYINPUT79), .B2(G169gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT81), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(G169gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(G176gat), .B1(new_n406_), .B2(KEYINPUT80), .ZN(new_n407_));
  OR2_X1    g206(.A1(KEYINPUT79), .A2(G169gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(KEYINPUT79), .A2(G169gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(KEYINPUT22), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n407_), .A2(new_n410_), .A3(new_n411_), .A4(new_n401_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n390_), .A2(new_n392_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n375_), .A2(new_n370_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n405_), .A2(new_n388_), .A3(new_n412_), .A4(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n369_), .A2(new_n397_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT20), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n373_), .A2(G190gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n370_), .A2(KEYINPUT26), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n376_), .A2(new_n378_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n394_), .A2(KEYINPUT90), .A3(new_n395_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT90), .B1(new_n394_), .B2(new_n395_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n389_), .B(new_n423_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT91), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n394_), .A2(new_n428_), .A3(new_n415_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n416_), .A2(KEYINPUT91), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n385_), .A2(KEYINPUT22), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n406_), .A2(new_n432_), .A3(new_n386_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n388_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n347_), .A2(G197gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n350_), .A2(G204gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT21), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n364_), .A2(new_n438_), .A3(new_n356_), .A4(new_n358_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n361_), .A2(new_n362_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n353_), .A2(new_n359_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT92), .B1(new_n435_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n423_), .A2(new_n389_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n394_), .A2(new_n395_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n444_), .B1(new_n447_), .B2(new_n424_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n433_), .A2(new_n388_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n449_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n442_), .B(KEYINPUT92), .C1(new_n448_), .C2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n420_), .B1(new_n443_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n416_), .A2(new_n388_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n407_), .A2(new_n410_), .A3(new_n401_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(KEYINPUT81), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n457_), .A2(new_n412_), .B1(new_n384_), .B2(new_n396_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n454_), .B1(new_n458_), .B2(new_n369_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(new_n419_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n342_), .B(new_n346_), .C1(new_n453_), .C2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n346_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n448_), .A2(new_n450_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n454_), .B1(new_n463_), .B2(new_n369_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n397_), .A2(new_n417_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT94), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n442_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n465_), .B2(new_n442_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n462_), .B(new_n464_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n461_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n418_), .A2(KEYINPUT20), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT89), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n442_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT92), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n451_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n477_), .A3(new_n420_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n342_), .B1(new_n478_), .B2(new_n346_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n341_), .B1(new_n471_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n346_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT93), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n482_), .A2(new_n340_), .A3(new_n470_), .A4(new_n461_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT103), .B(KEYINPUT27), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT102), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n464_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n346_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n473_), .A2(new_n477_), .A3(new_n462_), .A4(new_n420_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n488_), .B1(new_n492_), .B2(new_n341_), .ZN(new_n493_));
  AOI211_X1 g292(.A(KEYINPUT102), .B(new_n340_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n483_), .B(KEYINPUT27), .C1(new_n493_), .C2(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n487_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G155gat), .A2(G162gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(KEYINPUT1), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT1), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n500_), .A2(KEYINPUT84), .A3(G155gat), .A4(G162gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(KEYINPUT1), .ZN(new_n502_));
  OR2_X1    g301(.A1(G155gat), .A2(G162gat), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n499_), .A2(new_n501_), .A3(new_n502_), .A4(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G141gat), .B(G148gat), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT3), .ZN(new_n507_));
  INV_X1    g306(.A(G141gat), .ZN(new_n508_));
  INV_X1    g307(.A(G148gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G141gat), .A2(G148gat), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT2), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n510_), .A2(new_n513_), .A3(new_n514_), .A4(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(new_n498_), .A3(new_n503_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n506_), .A2(new_n517_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(KEYINPUT29), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n519_), .A2(KEYINPUT28), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(KEYINPUT28), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n369_), .B1(KEYINPUT29), .B2(new_n518_), .ZN(new_n522_));
  OR3_X1    g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n522_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G228gat), .A2(G233gat), .ZN(new_n525_));
  INV_X1    g324(.A(G78gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(new_n240_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G22gat), .B(G50gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n523_), .A2(new_n524_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G1gat), .B(G29gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G85gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT0), .B(G57gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(G134gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G127gat), .ZN(new_n540_));
  INV_X1    g339(.A(G127gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(G134gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(G120gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(G113gat), .ZN(new_n545_));
  INV_X1    g344(.A(G113gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(G120gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT82), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n540_), .A2(new_n542_), .A3(new_n545_), .A4(new_n547_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n543_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n553_), .A2(KEYINPUT82), .A3(new_n545_), .A4(new_n547_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n518_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G225gat), .A2(G233gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(new_n551_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n506_), .A2(new_n517_), .A3(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n556_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT97), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT97), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n556_), .A2(new_n562_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n557_), .B(KEYINPUT96), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n554_), .A2(new_n552_), .B1(new_n506_), .B2(new_n517_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n559_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT4), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT4), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n556_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n566_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n538_), .B1(new_n564_), .B2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n570_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n567_), .A2(KEYINPUT4), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n565_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(new_n537_), .A3(new_n561_), .A4(new_n563_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(KEYINPUT100), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT100), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n579_), .B(new_n538_), .C1(new_n564_), .C2(new_n572_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT101), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(KEYINPUT101), .A3(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n555_), .B(KEYINPUT31), .Z(new_n587_));
  XNOR2_X1  g386(.A(G71gat), .B(G99gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G43gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n465_), .B(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G227gat), .A2(G233gat), .ZN(new_n591_));
  INV_X1    g390(.A(G15gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT30), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n590_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT83), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n587_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n597_), .B1(new_n596_), .B2(new_n595_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n595_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(KEYINPUT83), .A3(new_n587_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n586_), .A2(new_n601_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n496_), .A2(new_n533_), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n557_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n556_), .A2(new_n565_), .A3(new_n559_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n538_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n606_), .B1(new_n577_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n577_), .A2(new_n607_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n577_), .A2(KEYINPUT98), .A3(new_n607_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n608_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n613_), .A2(new_n480_), .A3(new_n483_), .A4(KEYINPUT99), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n340_), .A2(KEYINPUT32), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n581_), .B1(new_n492_), .B2(new_n618_), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n471_), .A2(new_n479_), .A3(new_n618_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n616_), .A2(new_n617_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n533_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n533_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n487_), .A2(new_n624_), .A3(new_n495_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT104), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n487_), .A2(new_n624_), .A3(new_n627_), .A4(new_n495_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(new_n626_), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n603_), .B1(new_n629_), .B2(new_n601_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT75), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n233_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(new_n321_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n632_), .A2(new_n321_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n256_), .A2(new_n321_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n634_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G113gat), .B(G141gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT76), .ZN(new_n642_));
  XOR2_X1   g441(.A(G169gat), .B(G197gat), .Z(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n640_), .B(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n335_), .A2(new_n630_), .A3(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n315_), .A3(new_n586_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT38), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n645_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n310_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n268_), .A2(new_n270_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR4_X1   g453(.A1(new_n630_), .A2(new_n652_), .A3(new_n333_), .A4(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n315_), .B1(new_n655_), .B2(new_n586_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n649_), .A2(new_n650_), .A3(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT105), .Z(G1324gat));
  INV_X1    g457(.A(new_n496_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n646_), .A2(new_n316_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n655_), .A2(new_n659_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n662_), .B2(G8gat), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT39), .B(new_n316_), .C1(new_n655_), .C2(new_n659_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g465(.A(new_n601_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n592_), .B1(new_n655_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT41), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n646_), .A2(new_n592_), .A3(new_n667_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  INV_X1    g471(.A(new_n533_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n646_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n655_), .A2(new_n673_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(G22gat), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT42), .B(new_n672_), .C1(new_n655_), .C2(new_n673_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT106), .Z(G1327gat));
  NAND2_X1  g479(.A1(new_n654_), .A2(new_n333_), .ZN(new_n681_));
  NOR4_X1   g480(.A1(new_n630_), .A2(new_n645_), .A3(new_n309_), .A4(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n586_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n652_), .A2(new_n334_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n626_), .A2(new_n628_), .ZN(new_n687_));
  AOI22_X1  g486(.A1(new_n614_), .A2(new_n615_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n673_), .B1(new_n688_), .B2(new_n617_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n601_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n603_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n273_), .A2(new_n274_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n686_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n630_), .A2(KEYINPUT43), .A3(new_n275_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n684_), .B(new_n685_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n685_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n692_), .A2(new_n686_), .A3(new_n693_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n630_), .B2(new_n275_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n701_));
  OAI21_X1  g500(.A(new_n696_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n586_), .A2(G29gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n683_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n682_), .A2(new_n706_), .A3(new_n659_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT45), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n706_), .B1(new_n702_), .B2(new_n659_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n700_), .A2(new_n701_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n496_), .B1(new_n712_), .B2(new_n696_), .ZN(new_n713_));
  OAI211_X1 g512(.A(KEYINPUT46), .B(new_n708_), .C1(new_n713_), .C2(new_n706_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(G1329gat));
  INV_X1    g514(.A(G43gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n682_), .A2(new_n716_), .A3(new_n667_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n601_), .B1(new_n712_), .B2(new_n696_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n717_), .B(new_n718_), .C1(new_n719_), .C2(new_n716_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n718_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n716_), .B1(new_n702_), .B2(new_n667_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n717_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n720_), .A2(new_n724_), .ZN(G1330gat));
  AOI21_X1  g524(.A(G50gat), .B1(new_n682_), .B2(new_n673_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n673_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n702_), .B2(new_n727_), .ZN(G1331gat));
  NOR2_X1   g527(.A1(new_n693_), .A2(new_n333_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n692_), .A2(new_n645_), .A3(new_n309_), .A4(new_n729_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT109), .Z(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT110), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(KEYINPUT110), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n586_), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G57gat), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n334_), .A2(new_n645_), .ZN(new_n736_));
  NOR4_X1   g535(.A1(new_n630_), .A2(new_n310_), .A3(new_n654_), .A4(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n585_), .A2(new_n735_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n734_), .A2(new_n735_), .B1(new_n737_), .B2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n737_), .B2(new_n659_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT48), .Z(new_n742_));
  NAND2_X1  g541(.A1(new_n659_), .A2(new_n740_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT111), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n731_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n742_), .A2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n737_), .B2(new_n667_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT49), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n731_), .A2(new_n747_), .A3(new_n667_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1334gat));
  AOI21_X1  g550(.A(new_n526_), .B1(new_n737_), .B2(new_n673_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT50), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n731_), .A2(new_n526_), .A3(new_n673_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n310_), .A2(new_n681_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n692_), .A2(new_n645_), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n692_), .A2(KEYINPUT112), .A3(new_n645_), .A4(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n221_), .A3(new_n586_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n698_), .A2(new_n699_), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n310_), .A2(new_n651_), .A3(new_n334_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n586_), .A3(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n762_), .B1(new_n768_), .B2(new_n221_), .ZN(G1336gat));
  NAND3_X1  g568(.A1(new_n761_), .A2(new_n222_), .A3(new_n659_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n766_), .A2(new_n659_), .A3(new_n767_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n222_), .ZN(G1337gat));
  NAND2_X1  g571(.A1(new_n667_), .A2(new_n241_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n667_), .B(new_n767_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(G99gat), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT51), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(G99gat), .ZN(new_n780_));
  INV_X1    g579(.A(new_n774_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n777_), .A3(KEYINPUT51), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n774_), .B(new_n783_), .C1(new_n775_), .C2(G99gat), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n778_), .A2(new_n782_), .A3(new_n784_), .ZN(G1338gat));
  NOR2_X1   g584(.A1(new_n533_), .A2(G106gat), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n761_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n761_), .A2(KEYINPUT116), .A3(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n767_), .A2(new_n673_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n793_));
  OR3_X1    g592(.A1(new_n793_), .A2(KEYINPUT52), .A3(new_n240_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT52), .B1(new_n793_), .B2(new_n240_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT53), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n791_), .A2(new_n796_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1339gat));
  OAI21_X1  g600(.A(KEYINPUT54), .B1(new_n335_), .B2(new_n651_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n729_), .A2(new_n803_), .A3(new_n645_), .A4(new_n310_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n303_), .B1(new_n297_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n295_), .A2(new_n289_), .A3(new_n296_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n809_), .A2(new_n297_), .A3(new_n806_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n805_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n298_), .A2(KEYINPUT55), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT56), .B(new_n807_), .C1(new_n813_), .C2(new_n809_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n812_), .A3(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT117), .B(new_n805_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n645_), .A2(new_n304_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n636_), .A2(new_n639_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n637_), .A2(new_n635_), .A3(new_n638_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n644_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n819_), .A2(new_n644_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT118), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n822_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n653_), .B1(new_n818_), .B2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI221_X1 g629(.A(new_n653_), .B1(KEYINPUT119), .B2(KEYINPUT57), .C1(new_n818_), .C2(new_n827_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n294_), .A2(new_n298_), .A3(new_n303_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n822_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n811_), .B2(new_n814_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n834_), .A2(KEYINPUT58), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(KEYINPUT58), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n693_), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n830_), .A2(new_n831_), .A3(new_n837_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n802_), .A2(new_n804_), .B1(new_n838_), .B2(new_n333_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n659_), .A2(new_n673_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n586_), .A3(new_n667_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n546_), .A3(new_n651_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n802_), .A2(new_n804_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n838_), .A2(new_n333_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n841_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(KEYINPUT59), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n645_), .B1(new_n845_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n843_), .B1(new_n851_), .B2(new_n546_), .ZN(G1340gat));
  OAI21_X1  g651(.A(new_n544_), .B1(new_n310_), .B2(KEYINPUT60), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n842_), .B(new_n853_), .C1(KEYINPUT60), .C2(new_n544_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n310_), .B1(new_n845_), .B2(new_n850_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n544_), .ZN(G1341gat));
  AOI21_X1  g655(.A(G127gat), .B1(new_n842_), .B2(new_n334_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n845_), .A2(new_n850_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n333_), .A2(KEYINPUT120), .ZN(new_n859_));
  MUX2_X1   g658(.A(KEYINPUT120), .B(new_n859_), .S(G127gat), .Z(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n858_), .B2(new_n860_), .ZN(G1342gat));
  NOR2_X1   g660(.A1(new_n275_), .A2(new_n539_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n842_), .A2(new_n654_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n539_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n862_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n845_), .B2(new_n850_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G134gat), .B1(new_n842_), .B2(new_n654_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT121), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n871_), .ZN(G1343gat));
  NAND4_X1  g671(.A1(new_n496_), .A2(new_n673_), .A3(new_n586_), .A4(new_n601_), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(KEYINPUT122), .Z(new_n874_));
  NAND2_X1  g673(.A1(new_n848_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n645_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT123), .B(G141gat), .Z(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1344gat));
  NOR2_X1   g677(.A1(new_n875_), .A2(new_n310_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n509_), .ZN(G1345gat));
  NOR2_X1   g679(.A1(new_n875_), .A2(new_n333_), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT61), .B(G155gat), .Z(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  INV_X1    g682(.A(new_n875_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G162gat), .B1(new_n884_), .B2(new_n654_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n693_), .A2(G162gat), .ZN(new_n886_));
  XOR2_X1   g685(.A(new_n886_), .B(KEYINPUT124), .Z(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n884_), .B2(new_n887_), .ZN(G1347gat));
  NOR4_X1   g687(.A1(new_n496_), .A2(new_n673_), .A3(new_n586_), .A4(new_n601_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n848_), .A2(new_n651_), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  OR3_X1    g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n385_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n890_), .B2(new_n385_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n406_), .A3(new_n432_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(G1348gat));
  AND2_X1   g694(.A1(new_n848_), .A2(new_n889_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n309_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n334_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n382_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n375_), .B2(new_n899_), .ZN(G1350gat));
  NAND4_X1  g700(.A1(new_n896_), .A2(new_n421_), .A3(new_n422_), .A4(new_n654_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n896_), .A2(new_n693_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n370_), .ZN(G1351gat));
  NAND2_X1  g703(.A1(new_n624_), .A2(new_n601_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n839_), .A2(new_n496_), .A3(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n651_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT125), .B(G197gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1352gat));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n309_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n910_), .B(new_n911_), .Z(G1353gat));
  AOI211_X1 g711(.A(KEYINPUT63), .B(G211gat), .C1(new_n906_), .C2(new_n334_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n906_), .A2(new_n334_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT63), .B(G211gat), .Z(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(G1354gat));
  NAND3_X1  g715(.A1(new_n906_), .A2(new_n355_), .A3(new_n654_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n906_), .A2(new_n693_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n355_), .ZN(G1355gat));
endmodule


