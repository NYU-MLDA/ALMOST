//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n570_, new_n571_, new_n572_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT19), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT89), .Z(new_n204_));
  XOR2_X1   g003(.A(G197gat), .B(G204gat), .Z(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT21), .B1(new_n205_), .B2(KEYINPUT87), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT87), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT21), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n211_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n211_), .A2(new_n209_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(KEYINPUT88), .A3(new_n205_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n212_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G183gat), .ZN(new_n222_));
  INV_X1    g021(.A(G190gat), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT23), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n225_), .B1(G183gat), .B2(G190gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n221_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT25), .B(G183gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT26), .B(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G169gat), .ZN(new_n233_));
  INV_X1    g032(.A(G176gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT24), .A3(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n235_), .A2(KEYINPUT24), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n232_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT23), .B1(new_n222_), .B2(new_n223_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(KEYINPUT81), .B(KEYINPUT23), .C1(new_n222_), .C2(new_n223_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n224_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n229_), .B1(new_n239_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT20), .B1(new_n219_), .B2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT88), .B1(new_n217_), .B2(new_n205_), .ZN(new_n247_));
  NOR4_X1   g046(.A1(new_n207_), .A2(new_n211_), .A3(new_n215_), .A4(new_n209_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n221_), .B1(new_n244_), .B2(new_n228_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n227_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n251_), .A2(new_n237_), .A3(new_n238_), .A4(new_n232_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n249_), .A2(new_n212_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n204_), .B1(new_n246_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G8gat), .B(G36gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G64gat), .B(G92gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n219_), .B2(new_n245_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n249_), .A2(new_n252_), .A3(new_n250_), .A4(new_n212_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n203_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n254_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT95), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT95), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n254_), .A2(new_n263_), .A3(new_n266_), .A4(new_n259_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n259_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n246_), .A2(new_n253_), .A3(new_n204_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n203_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n265_), .A2(KEYINPUT27), .A3(new_n267_), .A4(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT96), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT27), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n254_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n259_), .B1(new_n254_), .B2(new_n263_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n272_), .A2(new_n273_), .A3(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n275_), .A2(new_n276_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(KEYINPUT96), .A3(new_n274_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G228gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(G78gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G106gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G22gat), .B(G50gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT86), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT2), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G155gat), .ZN(new_n296_));
  INV_X1    g095(.A(G162gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(KEYINPUT83), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(G155gat), .B2(G162gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n295_), .A2(new_n298_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(KEYINPUT1), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n298_), .A2(new_n303_), .A3(new_n300_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT84), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n301_), .A2(KEYINPUT1), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT84), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n298_), .A2(new_n303_), .A3(new_n300_), .A4(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT85), .ZN(new_n310_));
  INV_X1    g109(.A(new_n293_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(new_n291_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n310_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n302_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n315_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(KEYINPUT29), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n219_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT28), .B1(new_n315_), .B2(KEYINPUT29), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n319_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n288_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(new_n321_), .A3(new_n287_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n282_), .A2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G113gat), .B(G120gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n315_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n333_), .B(new_n302_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G1gat), .B(G29gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(G57gat), .B(G85gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n332_), .A2(KEYINPUT4), .A3(new_n334_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT91), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT91), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n332_), .A2(new_n345_), .A3(KEYINPUT4), .A4(new_n334_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n335_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n332_), .B2(KEYINPUT4), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n342_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n341_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n349_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n336_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G43gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n245_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(G15gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT30), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n361_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n366_), .A2(new_n367_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n331_), .B(KEYINPUT31), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(new_n367_), .A3(new_n370_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n328_), .A2(new_n358_), .A3(new_n374_), .ZN(new_n375_));
  AND4_X1   g174(.A1(new_n352_), .A2(new_n281_), .A3(new_n327_), .A4(new_n356_), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT93), .B(KEYINPUT33), .Z(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT94), .B1(new_n351_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT94), .ZN(new_n379_));
  INV_X1    g178(.A(new_n377_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n379_), .B(new_n380_), .C1(new_n354_), .C2(new_n342_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n351_), .A2(KEYINPUT33), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n332_), .A2(KEYINPUT4), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(new_n348_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n347_), .A2(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n332_), .A2(new_n334_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n341_), .B1(new_n386_), .B2(new_n348_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n279_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .A4(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n269_), .A2(new_n270_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n254_), .A2(new_n263_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n259_), .A2(KEYINPUT32), .ZN(new_n392_));
  MUX2_X1   g191(.A(new_n390_), .B(new_n391_), .S(new_n392_), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n357_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n327_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n376_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n375_), .B1(new_n397_), .B2(new_n374_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G15gat), .B(G22gat), .ZN(new_n399_));
  INV_X1    g198(.A(G1gat), .ZN(new_n400_));
  INV_X1    g199(.A(G8gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT14), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G8gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  XNOR2_X1  g204(.A(G29gat), .B(G36gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G43gat), .B(G50gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT78), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n408_), .B(KEYINPUT15), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n410_), .B1(new_n405_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G229gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n405_), .A2(new_n408_), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n417_), .B(KEYINPUT79), .Z(new_n418_));
  AND2_X1   g217(.A1(new_n418_), .A2(new_n410_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n416_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G113gat), .B(G141gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G169gat), .B(G197gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n422_), .B(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n398_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G85gat), .B(G92gat), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G99gat), .A2(G106gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT6), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT7), .ZN(new_n432_));
  INV_X1    g231(.A(G99gat), .ZN(new_n433_));
  INV_X1    g232(.A(G106gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n437_), .B(KEYINPUT66), .Z(new_n438_));
  AOI21_X1  g237(.A(new_n429_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT8), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n439_), .B1(KEYINPUT67), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(KEYINPUT10), .B(G99gat), .Z(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n434_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT64), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n428_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n428_), .A2(KEYINPUT65), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT9), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n449_), .B(new_n450_), .C1(G85gat), .C2(G92gat), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n447_), .A2(new_n431_), .A3(new_n448_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n444_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G57gat), .B(G64gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT11), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT68), .ZN(new_n456_));
  XOR2_X1   g255(.A(G71gat), .B(G78gat), .Z(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(KEYINPUT11), .B2(new_n454_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n456_), .B(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n453_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n446_), .B(KEYINPUT64), .Z(new_n464_));
  NAND3_X1  g263(.A1(new_n451_), .A2(new_n431_), .A3(new_n448_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n452_), .A2(KEYINPUT70), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n444_), .A3(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n459_), .A2(new_n462_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G230gat), .A2(G233gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n466_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n475_), .B2(new_n459_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n463_), .A2(new_n472_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT69), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n453_), .B2(new_n460_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n475_), .A2(KEYINPUT69), .A3(new_n459_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n461_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n477_), .B1(new_n483_), .B2(new_n474_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G120gat), .B(G148gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT5), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G176gat), .B(G204gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n488_), .B(KEYINPUT71), .Z(new_n491_));
  OAI21_X1  g290(.A(new_n490_), .B1(new_n484_), .B2(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n492_), .A2(KEYINPUT13), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(KEYINPUT13), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G231gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n405_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(new_n459_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT17), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G127gat), .B(G155gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G183gat), .B(G211gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  OR3_X1    g304(.A1(new_n499_), .A2(new_n500_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(KEYINPUT17), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n499_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n470_), .A2(new_n411_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n475_), .B2(new_n408_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n514_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n511_), .B(new_n516_), .C1(new_n519_), .C2(new_n518_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT74), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT75), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G190gat), .B(G218gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G134gat), .B(G162gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT36), .Z(new_n529_));
  INV_X1    g328(.A(KEYINPUT74), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n521_), .A2(new_n522_), .A3(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n524_), .A2(new_n525_), .A3(new_n529_), .A4(new_n531_), .ZN(new_n532_));
  OR3_X1    g331(.A1(new_n523_), .A2(KEYINPUT36), .A3(new_n528_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n529_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(new_n523_), .B2(KEYINPUT74), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n525_), .B1(new_n536_), .B2(new_n531_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT76), .B(KEYINPUT37), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n529_), .B(KEYINPUT73), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n523_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n533_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT37), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n427_), .A2(new_n495_), .A3(new_n510_), .A4(new_n545_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n546_), .A2(G1gat), .A3(new_n358_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT97), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(KEYINPUT38), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(KEYINPUT38), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n538_), .A2(KEYINPUT98), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT98), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n552_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n555_), .A2(new_n398_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n495_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n426_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n509_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n400_), .B1(new_n560_), .B2(new_n357_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT99), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n549_), .A2(new_n550_), .A3(new_n562_), .ZN(G1324gat));
  AOI21_X1  g362(.A(new_n401_), .B1(new_n560_), .B2(new_n282_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT39), .Z(new_n565_));
  INV_X1    g364(.A(new_n546_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(new_n401_), .A3(new_n282_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g368(.A(new_n363_), .B1(new_n560_), .B2(new_n374_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT41), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n566_), .A2(new_n363_), .A3(new_n374_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(G1326gat));
  INV_X1    g372(.A(G22gat), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n560_), .B2(new_n327_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT42), .Z(new_n576_));
  NAND3_X1  g375(.A1(new_n566_), .A2(new_n574_), .A3(new_n327_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(G1327gat));
  NOR2_X1   g377(.A1(new_n555_), .A2(new_n510_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n579_), .A2(new_n427_), .A3(new_n495_), .ZN(new_n580_));
  INV_X1    g379(.A(G29gat), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n357_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT43), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n538_), .A2(new_n539_), .B1(KEYINPUT37), .B2(new_n543_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n395_), .A2(new_n396_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n376_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n374_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n375_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n583_), .B(new_n584_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT100), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n398_), .A2(KEYINPUT100), .A3(new_n583_), .A4(new_n584_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n398_), .A2(new_n584_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT43), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n591_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n557_), .A2(new_n558_), .A3(new_n510_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT44), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n595_), .A2(KEYINPUT44), .A3(new_n596_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n600_), .A2(new_n358_), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n582_), .B1(new_n603_), .B2(new_n581_), .ZN(G1328gat));
  INV_X1    g403(.A(G36gat), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n580_), .A2(new_n605_), .A3(new_n282_), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT102), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n599_), .A2(KEYINPUT101), .A3(new_n282_), .A4(new_n601_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(G36gat), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n599_), .A2(new_n282_), .A3(new_n601_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT101), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n609_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n615_));
  AND4_X1   g414(.A1(new_n609_), .A2(new_n614_), .A3(G36gat), .A4(new_n610_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n608_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT46), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(KEYINPUT46), .B(new_n608_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1329gat));
  INV_X1    g420(.A(G43gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n580_), .A2(new_n622_), .A3(new_n374_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n600_), .A2(new_n373_), .A3(new_n602_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n624_), .B2(new_n622_), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(G1330gat));
  AOI21_X1  g426(.A(G50gat), .B1(new_n580_), .B2(new_n327_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n600_), .A2(new_n602_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n327_), .A2(G50gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n628_), .B1(new_n629_), .B2(new_n630_), .ZN(G1331gat));
  NOR2_X1   g430(.A1(new_n495_), .A2(new_n426_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n556_), .A2(new_n510_), .A3(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G57gat), .B1(new_n633_), .B2(new_n358_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n632_), .A2(new_n398_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n510_), .A3(new_n545_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT105), .Z(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n358_), .A2(G57gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n634_), .B1(new_n638_), .B2(new_n639_), .ZN(G1332gat));
  OAI21_X1  g439(.A(G64gat), .B1(new_n633_), .B2(new_n281_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT48), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n281_), .A2(G64gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n642_), .B1(new_n638_), .B2(new_n643_), .ZN(G1333gat));
  OAI21_X1  g443(.A(G71gat), .B1(new_n633_), .B2(new_n373_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT49), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n373_), .A2(G71gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n638_), .B2(new_n647_), .ZN(G1334gat));
  OAI21_X1  g447(.A(G78gat), .B1(new_n633_), .B2(new_n396_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT50), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n396_), .A2(G78gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(new_n638_), .B2(new_n651_), .ZN(G1335gat));
  NAND2_X1  g451(.A1(new_n635_), .A2(new_n579_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G85gat), .B1(new_n654_), .B2(new_n357_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT106), .Z(new_n656_));
  AND3_X1   g455(.A1(new_n595_), .A2(new_n509_), .A3(new_n632_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n357_), .A2(G85gat), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT107), .Z(new_n659_));
  AOI21_X1  g458(.A(new_n656_), .B1(new_n657_), .B2(new_n659_), .ZN(G1336gat));
  NOR3_X1   g459(.A1(new_n653_), .A2(G92gat), .A3(new_n281_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n282_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n662_), .B2(G92gat), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT108), .ZN(G1337gat));
  NAND3_X1  g463(.A1(new_n654_), .A2(new_n374_), .A3(new_n445_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n657_), .A2(new_n374_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n433_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g467(.A1(new_n654_), .A2(new_n434_), .A3(new_n327_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n595_), .A2(new_n327_), .A3(new_n509_), .A4(new_n632_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G106gat), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT109), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT52), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(KEYINPUT109), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n669_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g477(.A1(new_n545_), .A2(new_n495_), .A3(new_n558_), .A4(new_n510_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n679_), .B(new_n680_), .Z(new_n681_));
  AND2_X1   g480(.A1(new_n413_), .A2(new_n415_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n683_));
  MUX2_X1   g482(.A(new_n683_), .B(new_n420_), .S(new_n425_), .Z(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(new_n490_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n491_), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n461_), .A2(new_n462_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(KEYINPUT55), .A3(new_n476_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT113), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n477_), .A2(KEYINPUT113), .A3(KEYINPUT55), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n477_), .A2(KEYINPUT111), .A3(KEYINPUT55), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n687_), .A2(new_n476_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT55), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n690_), .B(new_n691_), .C1(new_n692_), .C2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT112), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n482_), .A2(new_n687_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n463_), .A2(new_n472_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT112), .B1(new_n700_), .B2(new_n481_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n473_), .B1(new_n699_), .B2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT56), .B(new_n686_), .C1(new_n697_), .C2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n699_), .A2(new_n701_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n474_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT111), .B1(new_n477_), .B2(KEYINPUT55), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n694_), .A2(new_n693_), .A3(new_n695_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n705_), .A2(new_n708_), .A3(new_n690_), .A4(new_n691_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT56), .B1(new_n709_), .B2(new_n686_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n703_), .B1(new_n710_), .B2(KEYINPUT117), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n686_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT56), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n712_), .A2(KEYINPUT117), .A3(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n685_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT58), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n545_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(KEYINPUT58), .B(new_n685_), .C1(new_n711_), .C2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n712_), .A2(KEYINPUT114), .A3(new_n713_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n426_), .A2(new_n490_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n703_), .A2(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n720_), .B(new_n722_), .C1(new_n724_), .C2(new_n710_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT115), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n492_), .B2(new_n684_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n492_), .A2(new_n726_), .A3(new_n684_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n554_), .B1(new_n725_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT57), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT57), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n728_), .A2(new_n729_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n724_), .A2(new_n710_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n721_), .B1(new_n710_), .B2(KEYINPUT114), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n737_), .B2(new_n554_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n719_), .A2(new_n732_), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n681_), .B1(new_n739_), .B2(new_n509_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n328_), .A2(new_n357_), .A3(new_n374_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n741_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n738_), .B(KEYINPUT116), .ZN(new_n746_));
  AOI22_X1  g545(.A1(new_n717_), .A2(new_n718_), .B1(KEYINPUT57), .B2(new_n731_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n681_), .B1(new_n748_), .B2(new_n509_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n742_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT59), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n745_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G113gat), .B1(new_n752_), .B2(new_n558_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n748_), .A2(new_n509_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n681_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n743_), .ZN(new_n757_));
  OR3_X1    g556(.A1(new_n757_), .A2(G113gat), .A3(new_n558_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n753_), .A2(new_n758_), .ZN(G1340gat));
  OAI21_X1  g558(.A(G120gat), .B1(new_n752_), .B2(new_n495_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT60), .ZN(new_n761_));
  AOI21_X1  g560(.A(G120gat), .B1(new_n557_), .B2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n761_), .B2(G120gat), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT119), .B1(new_n757_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n750_), .A2(new_n766_), .A3(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n760_), .A2(new_n768_), .ZN(G1341gat));
  OAI21_X1  g568(.A(G127gat), .B1(new_n752_), .B2(new_n509_), .ZN(new_n770_));
  OR3_X1    g569(.A1(new_n757_), .A2(G127gat), .A3(new_n509_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1342gat));
  INV_X1    g571(.A(KEYINPUT120), .ZN(new_n773_));
  INV_X1    g572(.A(G134gat), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n773_), .B(new_n774_), .C1(new_n757_), .C2(new_n555_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n749_), .A2(new_n555_), .A3(new_n742_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT120), .B1(new_n776_), .B2(G134gat), .ZN(new_n777_));
  INV_X1    g576(.A(new_n745_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n757_), .B2(KEYINPUT59), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n545_), .A2(new_n774_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n775_), .A2(new_n777_), .B1(new_n779_), .B2(new_n780_), .ZN(G1343gat));
  XNOR2_X1  g580(.A(KEYINPUT121), .B(G141gat), .ZN(new_n782_));
  NOR4_X1   g581(.A1(new_n374_), .A2(new_n358_), .A3(new_n282_), .A4(new_n396_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n756_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n782_), .B1(new_n785_), .B2(new_n426_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n782_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n784_), .A2(new_n558_), .A3(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1344gat));
  OR3_X1    g588(.A1(new_n784_), .A2(G148gat), .A3(new_n495_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G148gat), .B1(new_n784_), .B2(new_n495_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1345gat));
  XNOR2_X1  g591(.A(KEYINPUT61), .B(G155gat), .ZN(new_n793_));
  OR3_X1    g592(.A1(new_n784_), .A2(new_n509_), .A3(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n784_), .B2(new_n509_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1346gat));
  OAI21_X1  g595(.A(G162gat), .B1(new_n784_), .B2(new_n545_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n554_), .A2(new_n297_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n784_), .B2(new_n798_), .ZN(G1347gat));
  INV_X1    g598(.A(KEYINPUT124), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n357_), .A2(new_n373_), .A3(new_n281_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n327_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n510_), .B1(new_n747_), .B2(new_n738_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n426_), .B(new_n803_), .C1(new_n804_), .C2(new_n681_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n805_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT123), .B1(new_n805_), .B2(G169gat), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT123), .ZN(new_n810_));
  INV_X1    g609(.A(new_n803_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n740_), .A2(new_n558_), .A3(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n810_), .B(new_n808_), .C1(new_n812_), .C2(new_n233_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT22), .B(G169gat), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n800_), .B1(new_n809_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n810_), .B1(new_n812_), .B2(new_n233_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n805_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n819_));
  INV_X1    g618(.A(new_n808_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n821_), .A2(KEYINPUT124), .A3(new_n813_), .A4(new_n815_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n822_), .ZN(G1348gat));
  NOR2_X1   g622(.A1(new_n740_), .A2(new_n811_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G176gat), .B1(new_n824_), .B2(new_n557_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n749_), .A2(new_n327_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n495_), .A2(new_n234_), .A3(new_n802_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(G1349gat));
  NOR2_X1   g627(.A1(new_n802_), .A2(new_n509_), .ZN(new_n829_));
  AOI21_X1  g628(.A(G183gat), .B1(new_n826_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT125), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n509_), .A2(new_n230_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n824_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n831_), .B1(new_n824_), .B2(new_n832_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n830_), .A2(new_n833_), .A3(new_n834_), .ZN(G1350gat));
  NAND3_X1  g634(.A1(new_n824_), .A2(new_n231_), .A3(new_n554_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n740_), .A2(new_n545_), .A3(new_n811_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n223_), .ZN(G1351gat));
  NOR4_X1   g637(.A1(new_n374_), .A2(new_n396_), .A3(new_n357_), .A4(new_n281_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n749_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n426_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n557_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n510_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT63), .B(G211gat), .Z(new_n849_));
  NAND4_X1  g648(.A1(new_n756_), .A2(new_n510_), .A3(new_n839_), .A4(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT126), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT126), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n841_), .A2(new_n852_), .A3(new_n510_), .A4(new_n849_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n848_), .A2(new_n851_), .A3(new_n853_), .ZN(G1354gat));
  AOI21_X1  g653(.A(G218gat), .B1(new_n841_), .B2(new_n554_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n584_), .A2(G218gat), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT127), .Z(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n841_), .B2(new_n857_), .ZN(G1355gat));
endmodule


