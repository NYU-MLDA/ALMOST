//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n562_, new_n563_,
    new_n564_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT24), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  MUX2_X1   g003(.A(new_n203_), .B(KEYINPUT24), .S(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT23), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT25), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT80), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(KEYINPUT25), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n205_), .B(new_n207_), .C1(new_n210_), .C2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(new_n206_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(new_n216_), .B2(new_n206_), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT81), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT22), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n219_), .B(new_n222_), .C1(new_n223_), .C2(new_n220_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n218_), .A2(new_n224_), .A3(new_n202_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n214_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G227gat), .A2(G233gat), .ZN(new_n227_));
  INV_X1    g026(.A(G15gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT30), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n226_), .B(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G113gat), .B(G120gat), .Z(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT82), .B1(new_n234_), .B2(KEYINPUT31), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(KEYINPUT31), .B2(new_n234_), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n231_), .B(new_n236_), .Z(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G99gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G43gat), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(G141gat), .A2(G148gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G155gat), .A2(G162gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT83), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n248_));
  AND2_X1   g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(G155gat), .A3(G162gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT84), .Z(new_n252_));
  OAI211_X1 g051(.A(new_n244_), .B(new_n245_), .C1(new_n250_), .C2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n249_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT3), .B1(new_n245_), .B2(KEYINPUT85), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT2), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n244_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n245_), .A2(KEYINPUT85), .A3(KEYINPUT3), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n247_), .B(new_n254_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n253_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT29), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT89), .B(G204gat), .Z(new_n264_));
  OR3_X1    g063(.A1(new_n264_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n266_), .A2(KEYINPUT21), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n264_), .A2(G197gat), .ZN(new_n268_));
  INV_X1    g067(.A(G204gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT90), .B1(new_n269_), .B2(G197gat), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n265_), .B(new_n267_), .C1(new_n268_), .C2(new_n270_), .ZN(new_n271_));
  MUX2_X1   g070(.A(G204gat), .B(new_n264_), .S(G197gat), .Z(new_n272_));
  NAND2_X1  g071(.A1(KEYINPUT91), .A2(KEYINPUT21), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n266_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n263_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT88), .ZN(new_n278_));
  OAI21_X1  g077(.A(G233gat), .B1(new_n278_), .B2(G228gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n278_), .B2(G228gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT87), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n280_), .B1(new_n276_), .B2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n282_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G78gat), .B(G106gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n286_), .B(KEYINPUT93), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n284_), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n285_), .B(KEYINPUT92), .Z(new_n289_));
  AND2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n262_), .A2(KEYINPUT29), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G22gat), .B(G50gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  OR3_X1    g094(.A1(new_n287_), .A2(new_n290_), .A3(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n288_), .A2(new_n289_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n295_), .B1(new_n290_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G8gat), .B(G36gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  NAND2_X1  g103(.A1(new_n209_), .A2(new_n212_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n211_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(new_n205_), .A3(new_n207_), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT22), .B(G169gat), .Z(new_n309_));
  OAI211_X1 g108(.A(new_n218_), .B(new_n202_), .C1(G176gat), .C2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n276_), .A2(new_n311_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n312_), .B(KEYINPUT20), .C1(new_n276_), .C2(new_n226_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT19), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n276_), .A2(new_n226_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n317_), .B(KEYINPUT20), .C1(new_n276_), .C2(new_n311_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(new_n315_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n304_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT95), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n316_), .A2(new_n319_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n304_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n321_), .B(new_n324_), .Z(new_n325_));
  INV_X1    g124(.A(new_n234_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n326_), .B1(new_n253_), .B2(new_n261_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n262_), .A2(new_n234_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(new_n327_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n331_), .B2(KEYINPUT4), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n333_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G85gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT0), .B(G57gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT33), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT33), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n332_), .A2(new_n333_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n341_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n325_), .B(new_n344_), .C1(new_n343_), .C2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n343_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n337_), .A2(new_n342_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n323_), .A2(KEYINPUT32), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n322_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT96), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n313_), .A2(new_n315_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n318_), .A2(new_n315_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n352_), .B(new_n354_), .C1(new_n359_), .C2(new_n353_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n299_), .B1(new_n349_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT97), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n325_), .A2(KEYINPUT27), .ZN(new_n363_));
  OAI211_X1 g162(.A(KEYINPUT27), .B(new_n324_), .C1(new_n359_), .C2(new_n323_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n352_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n299_), .A2(new_n366_), .ZN(new_n367_));
  OAI22_X1  g166(.A1(new_n361_), .A2(new_n362_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  AOI211_X1 g167(.A(KEYINPUT97), .B(new_n299_), .C1(new_n360_), .C2(new_n349_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n243_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n365_), .A2(new_n299_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n352_), .A2(new_n243_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G15gat), .B(G22gat), .Z(new_n375_));
  NAND2_X1  g174(.A1(G1gat), .A2(G8gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(KEYINPUT14), .B2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT78), .ZN(new_n378_));
  XOR2_X1   g177(.A(G1gat), .B(G8gat), .Z(new_n379_));
  AND2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n378_), .A2(new_n379_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G29gat), .B(G36gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT74), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G43gat), .B(G50gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n378_), .B(new_n379_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n386_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G229gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n386_), .B(KEYINPUT15), .Z(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n389_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n388_), .A3(new_n392_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G113gat), .B(G141gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT79), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G169gat), .B(G197gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n400_), .B(new_n401_), .Z(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n394_), .A2(new_n397_), .A3(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n374_), .A2(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(G230gat), .A2(G233gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(G99gat), .A2(G106gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT7), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(KEYINPUT65), .B2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(KEYINPUT65), .B(KEYINPUT7), .Z(new_n413_));
  AOI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(new_n410_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G99gat), .A2(G106gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT6), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT8), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G85gat), .B(G92gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT67), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT66), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT66), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT6), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n424_), .A2(new_n426_), .A3(new_n415_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n415_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n422_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n415_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n425_), .A2(KEYINPUT6), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n423_), .A2(KEYINPUT66), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n424_), .A2(new_n426_), .A3(new_n415_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(KEYINPUT67), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n429_), .A2(new_n435_), .A3(new_n414_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT68), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n420_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT8), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n436_), .B2(new_n420_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n421_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G57gat), .B(G64gat), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n444_));
  XOR2_X1   g243(.A(G71gat), .B(G78gat), .Z(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n444_), .A2(new_n445_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT9), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(G85gat), .A3(G92gat), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n416_), .B(new_n450_), .C1(new_n449_), .C2(new_n419_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT10), .B(G99gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n452_), .B(KEYINPUT64), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G106gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n451_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n441_), .A2(new_n448_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n436_), .A2(new_n420_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT68), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(KEYINPUT8), .A3(new_n438_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n456_), .B1(new_n463_), .B2(new_n421_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(KEYINPUT69), .A3(new_n448_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n464_), .A2(new_n448_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n409_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n464_), .B2(new_n448_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n409_), .B1(new_n464_), .B2(new_n448_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n441_), .A2(KEYINPUT70), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT70), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n473_), .B(new_n421_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n456_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n446_), .A2(KEYINPUT12), .A3(new_n447_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n470_), .B(new_n471_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G120gat), .B(G148gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT5), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G176gat), .B(G204gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n468_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT72), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n468_), .A2(KEYINPUT72), .A3(new_n477_), .A4(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n468_), .A2(new_n477_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n481_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(KEYINPUT13), .A3(new_n489_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n495_), .A2(KEYINPUT73), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(KEYINPUT73), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n448_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n389_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G127gat), .B(G155gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT16), .ZN(new_n505_));
  XOR2_X1   g304(.A(G183gat), .B(G211gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n502_), .A2(new_n503_), .A3(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(KEYINPUT17), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n502_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT35), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT34), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n464_), .A2(new_n387_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n395_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n516_), .B1(new_n475_), .B2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n515_), .A2(new_n512_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI221_X1 g319(.A(new_n516_), .B1(new_n512_), .B2(new_n515_), .C1(new_n475_), .C2(new_n517_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G190gat), .B(G218gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT75), .ZN(new_n523_));
  XOR2_X1   g322(.A(G134gat), .B(G162gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(KEYINPUT36), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n520_), .A2(new_n521_), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT76), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT76), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n520_), .A2(new_n521_), .A3(new_n530_), .A4(new_n527_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n525_), .B(KEYINPUT36), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT77), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT37), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NOR4_X1   g341(.A1(new_n408_), .A2(new_n499_), .A3(new_n511_), .A4(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(G1gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n352_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT38), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n532_), .A2(new_n536_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n494_), .A2(new_n406_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n550_), .A2(new_n510_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n544_), .B1(new_n552_), .B2(new_n352_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n546_), .B2(new_n545_), .ZN(G1324gat));
  INV_X1    g354(.A(G8gat), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n552_), .B2(new_n365_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT39), .Z(new_n558_));
  NAND3_X1  g357(.A1(new_n543_), .A2(new_n556_), .A3(new_n365_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n560_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g360(.A(new_n228_), .B1(new_n552_), .B2(new_n242_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT41), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n543_), .A2(new_n228_), .A3(new_n242_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(G1326gat));
  INV_X1    g364(.A(G22gat), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n552_), .B2(new_n299_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT42), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n299_), .A2(new_n566_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT98), .Z(new_n570_));
  NAND2_X1  g369(.A1(new_n543_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(G1327gat));
  INV_X1    g371(.A(KEYINPUT101), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n548_), .A2(new_n510_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n495_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n408_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n374_), .A2(KEYINPUT101), .A3(new_n407_), .A4(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(G29gat), .B1(new_n579_), .B2(new_n352_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n374_), .A2(new_n542_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT43), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT100), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n542_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n374_), .B(new_n542_), .C1(new_n583_), .C2(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n551_), .A2(new_n511_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT99), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT44), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n352_), .A2(G29gat), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n580_), .B1(new_n591_), .B2(new_n592_), .ZN(G1328gat));
  XOR2_X1   g392(.A(new_n590_), .B(KEYINPUT44), .Z(new_n594_));
  INV_X1    g393(.A(new_n365_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G36gat), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(G36gat), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n576_), .A2(new_n578_), .A3(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT45), .Z(new_n600_));
  NOR2_X1   g399(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n596_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n597_), .B1(new_n596_), .B2(new_n602_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(G1329gat));
  AOI21_X1  g404(.A(G43gat), .B1(new_n579_), .B2(new_n242_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n242_), .A2(G43gat), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n591_), .B2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(G1330gat));
  INV_X1    g409(.A(new_n299_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G50gat), .B1(new_n594_), .B2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(G50gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT104), .Z(new_n614_));
  NAND2_X1  g413(.A1(new_n579_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(G1331gat));
  AOI21_X1  g415(.A(new_n407_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n538_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n548_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n539_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n617_), .A2(new_n494_), .A3(new_n510_), .A4(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT105), .Z(new_n622_));
  INV_X1    g421(.A(G57gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n352_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n407_), .A2(new_n511_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n550_), .A2(new_n499_), .A3(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G57gat), .B1(new_n626_), .B2(new_n366_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(G1332gat));
  INV_X1    g427(.A(G64gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n622_), .A2(new_n629_), .A3(new_n365_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G64gat), .B1(new_n626_), .B2(new_n595_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT48), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(G1333gat));
  INV_X1    g432(.A(G71gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n622_), .A2(new_n634_), .A3(new_n242_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G71gat), .B1(new_n626_), .B2(new_n243_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT49), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1334gat));
  INV_X1    g437(.A(G78gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n622_), .A2(new_n639_), .A3(new_n299_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G78gat), .B1(new_n626_), .B2(new_n611_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT50), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(G1335gat));
  AND2_X1   g442(.A1(new_n617_), .A2(new_n574_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n499_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G85gat), .B1(new_n646_), .B2(new_n352_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n495_), .A2(new_n407_), .A3(new_n510_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n352_), .A2(G85gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT106), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n647_), .B1(new_n650_), .B2(new_n652_), .ZN(G1336gat));
  AOI21_X1  g452(.A(G92gat), .B1(new_n646_), .B2(new_n365_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT107), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n365_), .A2(G92gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT108), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n650_), .B2(new_n657_), .ZN(G1337gat));
  INV_X1    g457(.A(KEYINPUT110), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n646_), .A2(new_n454_), .A3(new_n242_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n650_), .A2(new_n242_), .ZN(new_n661_));
  INV_X1    g460(.A(G99gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n660_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n663_), .B2(KEYINPUT51), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(KEYINPUT109), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT51), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n663_), .B2(KEYINPUT109), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n664_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n665_), .A2(new_n667_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(KEYINPUT110), .B2(new_n669_), .ZN(G1338gat));
  NAND3_X1  g469(.A1(new_n646_), .A2(new_n455_), .A3(new_n299_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT52), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT111), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n650_), .A2(new_n673_), .A3(new_n299_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(G106gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n650_), .A2(new_n299_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT111), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n672_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  AND4_X1   g477(.A1(new_n672_), .A2(new_n677_), .A3(G106gat), .A4(new_n674_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n671_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT53), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT53), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n671_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1339gat));
  OAI21_X1  g483(.A(new_n470_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n409_), .B1(new_n685_), .B2(new_n466_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n474_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n473_), .B1(new_n463_), .B2(new_n421_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n457_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n476_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n691_), .A2(KEYINPUT55), .A3(new_n470_), .A4(new_n471_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT55), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n477_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n686_), .A2(new_n692_), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n481_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT56), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(KEYINPUT56), .A3(new_n481_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n404_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT113), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n396_), .A2(new_n388_), .A3(new_n393_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n701_), .B2(KEYINPUT113), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n405_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT58), .B1(new_n700_), .B2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT114), .B1(new_n620_), .B2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n700_), .A2(KEYINPUT58), .A3(new_n706_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n695_), .A2(KEYINPUT56), .A3(new_n481_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT56), .B1(new_n695_), .B2(new_n481_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n706_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT58), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT114), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n542_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n708_), .A2(new_n709_), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n705_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n490_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n406_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n720_));
  OAI22_X1  g519(.A1(KEYINPUT112), .A2(new_n720_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(KEYINPUT112), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n548_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT57), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(KEYINPUT57), .A3(new_n548_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n717_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n511_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n495_), .A2(new_n620_), .A3(new_n625_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(KEYINPUT54), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(KEYINPUT54), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n729_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n371_), .A2(new_n352_), .A3(new_n242_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT115), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(G113gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n407_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT117), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n717_), .A2(KEYINPUT116), .A3(new_n726_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT116), .B1(new_n717_), .B2(new_n726_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n727_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n746_), .B2(new_n510_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n717_), .A2(new_n726_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n717_), .A2(KEYINPUT116), .A3(new_n726_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(KEYINPUT117), .A3(new_n511_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n747_), .A2(new_n733_), .A3(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n735_), .A2(KEYINPUT59), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n728_), .A2(new_n511_), .B1(new_n732_), .B2(new_n731_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT59), .B1(new_n757_), .B2(new_n735_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(new_n407_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n741_), .B1(new_n760_), .B2(new_n740_), .ZN(G1340gat));
  INV_X1    g560(.A(G120gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n495_), .B2(KEYINPUT60), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n739_), .B(new_n763_), .C1(KEYINPUT60), .C2(new_n762_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n758_), .A2(new_n499_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G120gat), .B1(new_n766_), .B2(KEYINPUT118), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n768_), .B(new_n765_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT119), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT119), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n764_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1341gat));
  AOI21_X1  g573(.A(G127gat), .B1(new_n739_), .B2(new_n510_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n510_), .A2(G127gat), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT120), .Z(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n759_), .B2(new_n777_), .ZN(G1342gat));
  NAND3_X1  g577(.A1(new_n756_), .A2(new_n542_), .A3(new_n758_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(G134gat), .ZN(new_n780_));
  OR3_X1    g579(.A1(new_n738_), .A2(G134gat), .A3(new_n548_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT121), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n780_), .A2(new_n781_), .A3(KEYINPUT121), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1343gat));
  NOR2_X1   g585(.A1(new_n757_), .A2(new_n242_), .ZN(new_n787_));
  AND4_X1   g586(.A1(new_n299_), .A2(new_n787_), .A3(new_n352_), .A4(new_n595_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n407_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n499_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g591(.A1(new_n788_), .A2(new_n510_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT122), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT61), .B(G155gat), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n794_), .B(new_n796_), .ZN(G1346gat));
  INV_X1    g596(.A(G162gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n788_), .A2(new_n798_), .A3(new_n549_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n788_), .A2(new_n542_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n798_), .ZN(G1347gat));
  NAND2_X1  g600(.A1(new_n365_), .A2(new_n372_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n407_), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(KEYINPUT123), .Z(new_n805_));
  AOI21_X1  g604(.A(new_n510_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n733_), .B1(new_n806_), .B2(KEYINPUT117), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n746_), .A2(new_n742_), .A3(new_n510_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n611_), .B(new_n805_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT124), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G169gat), .B1(new_n809_), .B2(KEYINPUT124), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT62), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n809_), .A2(KEYINPUT124), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT62), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(G169gat), .A4(new_n810_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n754_), .A2(new_n611_), .ZN(new_n818_));
  OR3_X1    g617(.A1(new_n818_), .A2(new_n309_), .A3(new_n804_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1348gat));
  OAI211_X1 g619(.A(new_n611_), .B(new_n803_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(G176gat), .B1(new_n822_), .B2(new_n494_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n757_), .A2(new_n299_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n498_), .A2(new_n219_), .A3(new_n802_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(G1349gat));
  NAND2_X1  g625(.A1(new_n803_), .A2(new_n510_), .ZN(new_n827_));
  OR3_X1    g626(.A1(new_n818_), .A2(new_n306_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n824_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n208_), .B1(new_n829_), .B2(new_n827_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1350gat));
  OAI21_X1  g630(.A(G190gat), .B1(new_n821_), .B2(new_n620_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n549_), .A2(new_n211_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT125), .Z(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n821_), .B2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT126), .ZN(G1351gat));
  NOR2_X1   g635(.A1(new_n595_), .A2(new_n367_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n787_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n407_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g640(.A1(new_n838_), .A2(new_n498_), .ZN(new_n842_));
  MUX2_X1   g641(.A(G204gat), .B(new_n264_), .S(new_n842_), .Z(G1353gat));
  NOR2_X1   g642(.A1(new_n838_), .A2(new_n511_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n845_));
  AND2_X1   g644(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n844_), .B2(new_n845_), .ZN(G1354gat));
  AND3_X1   g647(.A1(new_n839_), .A2(G218gat), .A3(new_n542_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n838_), .A2(new_n548_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n850_), .A2(KEYINPUT127), .ZN(new_n851_));
  AOI21_X1  g650(.A(G218gat), .B1(new_n850_), .B2(KEYINPUT127), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n849_), .B1(new_n851_), .B2(new_n852_), .ZN(G1355gat));
endmodule


