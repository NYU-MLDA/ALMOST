//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT86), .ZN(new_n203_));
  INV_X1    g002(.A(G204gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n203_), .B1(new_n204_), .B2(G197gat), .ZN(new_n205_));
  INV_X1    g004(.A(G197gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n204_), .A2(G197gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT85), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n206_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(KEYINPUT87), .A2(KEYINPUT21), .ZN(new_n212_));
  NOR2_X1   g011(.A1(KEYINPUT87), .A2(KEYINPUT21), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .A4(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G218gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G211gat), .ZN(new_n217_));
  INV_X1    g016(.A(G211gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G218gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n206_), .A2(G204gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n209_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(KEYINPUT21), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n215_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n220_), .A2(KEYINPUT21), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT84), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G228gat), .A2(G233gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G155gat), .ZN(new_n232_));
  INV_X1    g031(.A(G162gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G155gat), .A3(G162gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR3_X1   g037(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n234_), .B(new_n236_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT82), .ZN(new_n241_));
  INV_X1    g040(.A(G141gat), .ZN(new_n242_));
  INV_X1    g041(.A(G148gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n244_), .A2(new_n245_), .B1(G141gat), .B2(G148gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n240_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT2), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n249_), .A2(new_n251_), .A3(new_n252_), .A4(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n256_), .A2(new_n237_), .B1(G155gat), .B2(G162gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n247_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT28), .B1(new_n259_), .B2(KEYINPUT29), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n240_), .A2(new_n246_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n231_), .A2(new_n260_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n264_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(new_n230_), .A3(new_n229_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n261_), .A2(new_n263_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n215_), .A2(new_n223_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n270_));
  OAI21_X1  g069(.A(G78gat), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n259_), .A2(KEYINPUT29), .ZN(new_n272_));
  INV_X1    g071(.A(G78gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n228_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n271_), .A2(new_n274_), .A3(G106gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(G106gat), .B1(new_n271_), .B2(new_n274_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G22gat), .B(G50gat), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n271_), .A2(new_n274_), .ZN(new_n281_));
  INV_X1    g080(.A(G106gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n280_), .B1(new_n283_), .B2(new_n275_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n268_), .B1(new_n279_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n278_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n275_), .A3(new_n280_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(new_n267_), .A4(new_n265_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT19), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT23), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(G183gat), .A3(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(G183gat), .B2(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT22), .B(G169gat), .ZN(new_n300_));
  INV_X1    g099(.A(G176gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G183gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT25), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT25), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G183gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT88), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT88), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n305_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT26), .B(G190gat), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n309_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n293_), .A2(new_n295_), .A3(KEYINPUT76), .ZN(new_n314_));
  INV_X1    g113(.A(G169gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n301_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(KEYINPUT24), .A3(new_n298_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT76), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n292_), .A2(new_n318_), .A3(KEYINPUT23), .ZN(new_n319_));
  OR3_X1    g118(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n314_), .A2(new_n317_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n303_), .B1(new_n313_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT20), .B1(new_n322_), .B2(new_n228_), .ZN(new_n323_));
  INV_X1    g122(.A(G190gat), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n305_), .B(new_n307_), .C1(KEYINPUT26), .C2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT73), .B1(new_n326_), .B2(G190gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(new_n324_), .A3(KEYINPUT26), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT74), .B1(new_n325_), .B2(new_n330_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n317_), .A2(new_n296_), .A3(new_n320_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n337_), .A2(new_n315_), .A3(KEYINPUT22), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(new_n315_), .B2(KEYINPUT22), .ZN(new_n339_));
  AOI21_X1  g138(.A(G176gat), .B1(new_n315_), .B2(KEYINPUT22), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n314_), .A2(new_n319_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  OAI221_X1 g142(.A(new_n298_), .B1(new_n338_), .B2(new_n341_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n270_), .B1(new_n336_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n291_), .B1(new_n323_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n347_));
  AND4_X1   g146(.A1(new_n319_), .A2(new_n314_), .A3(new_n317_), .A4(new_n320_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n309_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n348_), .A2(new_n349_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n347_), .B1(new_n350_), .B2(new_n270_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n322_), .A2(new_n228_), .A3(KEYINPUT89), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n336_), .A2(new_n344_), .A3(new_n270_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT20), .A4(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n346_), .B1(new_n354_), .B2(new_n291_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT18), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G64gat), .B(G92gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n291_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n359_), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n323_), .A2(new_n345_), .A3(new_n291_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(KEYINPUT27), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT94), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT27), .ZN(new_n367_));
  INV_X1    g166(.A(new_n364_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n362_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n367_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT94), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n360_), .A2(new_n364_), .A3(new_n371_), .A4(KEYINPUT27), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n289_), .A2(new_n366_), .A3(new_n370_), .A4(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT77), .B(KEYINPUT30), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n336_), .A2(new_n344_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n336_), .B2(new_n344_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT78), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n336_), .A2(new_n344_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n336_), .A2(new_n344_), .A3(new_n374_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G43gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(G15gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n385_), .B(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n377_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n388_), .ZN(new_n390_));
  OAI211_X1 g189(.A(KEYINPUT78), .B(new_n390_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n393_));
  XOR2_X1   g192(.A(G127gat), .B(G134gat), .Z(new_n394_));
  INV_X1    g193(.A(G120gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G113gat), .ZN(new_n396_));
  INV_X1    g195(.A(G113gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G120gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G127gat), .B(G134gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n393_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n394_), .A2(new_n399_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n402_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(KEYINPUT80), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(KEYINPUT81), .A3(new_n407_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(KEYINPUT31), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT79), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT31), .B1(new_n410_), .B2(new_n411_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n392_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n389_), .A2(new_n415_), .A3(new_n391_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G85gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT0), .B(G57gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n400_), .A2(new_n403_), .A3(new_n393_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT80), .B1(new_n405_), .B2(new_n406_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n259_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT90), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n247_), .B(new_n258_), .C1(new_n400_), .C2(new_n403_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n428_), .A2(KEYINPUT92), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n430_), .B(new_n431_), .C1(new_n408_), .C2(new_n261_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n427_), .A2(KEYINPUT91), .A3(new_n437_), .A4(new_n259_), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT4), .B(new_n431_), .C1(new_n408_), .C2(new_n261_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n259_), .A2(new_n404_), .A3(new_n437_), .A4(new_n407_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT91), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n430_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .A4(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n424_), .B1(new_n436_), .B2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n424_), .A3(new_n435_), .A4(new_n432_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT93), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n444_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n432_), .A2(new_n435_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n423_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT93), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n446_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n419_), .A2(new_n448_), .A3(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n202_), .B1(new_n373_), .B2(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n366_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n419_), .A2(new_n448_), .A3(new_n453_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n456_), .A2(KEYINPUT95), .A3(new_n289_), .A4(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .A4(new_n430_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n443_), .B(new_n431_), .C1(new_n408_), .C2(new_n261_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n460_), .A2(new_n423_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT33), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n446_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n361_), .A2(new_n363_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n359_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n436_), .A2(KEYINPUT33), .A3(new_n424_), .A4(new_n444_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n464_), .A2(new_n466_), .A3(new_n364_), .A4(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n355_), .A2(KEYINPUT32), .A3(new_n362_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n362_), .A2(KEYINPUT32), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n361_), .A2(new_n470_), .A3(new_n363_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n469_), .B(new_n471_), .C1(new_n445_), .C2(new_n447_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n289_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n366_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n448_), .A2(new_n453_), .A3(new_n288_), .A4(new_n285_), .ZN(new_n476_));
  OAI22_X1  g275(.A1(new_n473_), .A2(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n419_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n455_), .A2(new_n458_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G29gat), .B(G36gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G43gat), .B(G50gat), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G43gat), .B(G50gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  INV_X1    g288(.A(G1gat), .ZN(new_n490_));
  INV_X1    g289(.A(G8gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT14), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G1gat), .B(G8gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n483_), .A2(KEYINPUT15), .A3(new_n485_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n488_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n493_), .A2(new_n494_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n494_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n486_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n502_), .A2(KEYINPUT72), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n495_), .B(new_n486_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n502_), .B(KEYINPUT72), .C1(new_n504_), .C2(new_n498_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n503_), .A2(new_n505_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G120gat), .B(G148gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT5), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G176gat), .B(G204gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n519_));
  INV_X1    g318(.A(G99gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n282_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT65), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT6), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(KEYINPUT65), .ZN(new_n527_));
  OAI22_X1  g326(.A1(new_n525_), .A2(new_n527_), .B1(new_n520_), .B2(new_n282_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(KEYINPUT65), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(KEYINPUT6), .ZN(new_n530_));
  AND2_X1   g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n523_), .B1(new_n528_), .B2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G85gat), .B(G92gat), .Z(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT8), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT8), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n531_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n537_), .B(new_n534_), .C1(new_n540_), .C2(new_n523_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT66), .ZN(new_n543_));
  OR2_X1    g342(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n282_), .A3(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n547_));
  OAI211_X1 g346(.A(G85gat), .B(G92gat), .C1(KEYINPUT64), .C2(KEYINPUT9), .ZN(new_n548_));
  OAI211_X1 g347(.A(KEYINPUT64), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n543_), .B1(new_n547_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n528_), .A2(new_n532_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n555_), .A2(KEYINPUT66), .A3(new_n552_), .A4(new_n546_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n542_), .A2(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(G78gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n273_), .A3(new_n560_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G57gat), .B(G64gat), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n562_), .A2(new_n563_), .B1(KEYINPUT11), .B2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(KEYINPUT11), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n562_), .A2(new_n563_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n558_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n542_), .A2(new_n557_), .A3(new_n568_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(KEYINPUT68), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n568_), .B1(new_n542_), .B2(new_n557_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n572_), .A2(new_n574_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n570_), .A2(KEYINPUT12), .A3(new_n571_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT12), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n558_), .A2(new_n581_), .A3(new_n569_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n574_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n518_), .B1(new_n579_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n571_), .A2(KEYINPUT12), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(new_n575_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n582_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n573_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n518_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n578_), .A3(new_n589_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n584_), .A2(KEYINPUT13), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT13), .B1(new_n584_), .B2(new_n590_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT16), .ZN(new_n595_));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n495_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n568_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(new_n598_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n603_), .B2(new_n597_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT71), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n604_), .B(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT34), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n542_), .A2(new_n557_), .A3(new_n486_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n488_), .A2(new_n496_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n542_), .B2(new_n557_), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT35), .B(new_n609_), .C1(new_n610_), .C2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n611_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n558_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n542_), .A2(new_n557_), .A3(new_n486_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .A4(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT36), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT69), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT37), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n623_), .A2(KEYINPUT36), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n613_), .A2(new_n619_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT69), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n620_), .A2(new_n630_), .A3(new_n624_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n626_), .A2(new_n627_), .A3(new_n629_), .A4(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT70), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n625_), .A2(new_n629_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT37), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n632_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n633_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n593_), .B(new_n607_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n479_), .A2(new_n514_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n448_), .A2(new_n453_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n490_), .A3(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT96), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(KEYINPUT96), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT97), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT97), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT38), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n626_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT98), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n479_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n593_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n607_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n514_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n640_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n645_), .A2(KEYINPUT38), .A3(new_n646_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n649_), .A2(new_n659_), .A3(new_n660_), .ZN(G1324gat));
  NAND3_X1  g460(.A1(new_n639_), .A2(new_n491_), .A3(new_n475_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G8gat), .B1(new_n657_), .B2(new_n456_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n663_), .A2(KEYINPUT39), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(KEYINPUT39), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g466(.A(G15gat), .B1(new_n657_), .B2(new_n478_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT41), .Z(new_n669_));
  INV_X1    g468(.A(G15gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n639_), .A2(new_n670_), .A3(new_n419_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1326gat));
  XNOR2_X1  g471(.A(new_n289_), .B(KEYINPUT99), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G22gat), .B1(new_n657_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT42), .ZN(new_n676_));
  INV_X1    g475(.A(G22gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n639_), .A2(new_n677_), .A3(new_n673_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1327gat));
  INV_X1    g478(.A(new_n650_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n655_), .A2(new_n680_), .ZN(new_n681_));
  NOR4_X1   g480(.A1(new_n479_), .A2(new_n514_), .A3(new_n654_), .A4(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n640_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n655_), .A2(new_n513_), .A3(new_n593_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n632_), .A2(new_n635_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT70), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n632_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n479_), .A2(KEYINPUT43), .A3(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(KEYINPUT100), .B(KEYINPUT43), .Z(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n458_), .A2(new_n455_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n477_), .A2(new_n478_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n636_), .A2(new_n637_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT44), .B(new_n685_), .C1(new_n690_), .C2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT101), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n691_), .B1(new_n479_), .B2(new_n689_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n695_), .A2(new_n701_), .A3(new_n696_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n684_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n699_), .A2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n685_), .B1(new_n690_), .B2(new_n697_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n706_), .A2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n640_), .A2(G29gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n683_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  NOR2_X1   g511(.A1(new_n456_), .A2(G36gat), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n682_), .A2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(KEYINPUT45), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(KEYINPUT45), .ZN(new_n716_));
  OAI22_X1  g515(.A1(new_n715_), .A2(new_n716_), .B1(KEYINPUT102), .B2(KEYINPUT46), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n706_), .A2(new_n475_), .A3(new_n709_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G36gat), .ZN(new_n719_));
  AND2_X1   g518(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(G1329gat));
  NAND4_X1  g520(.A1(new_n706_), .A2(G43gat), .A3(new_n419_), .A4(new_n709_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G43gat), .B1(new_n682_), .B2(new_n419_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g525(.A(G50gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n673_), .A2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT105), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n682_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n474_), .B1(new_n703_), .B2(KEYINPUT44), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n699_), .B2(new_n705_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n727_), .B1(new_n732_), .B2(KEYINPUT103), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n289_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n706_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT104), .B1(new_n733_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n700_), .A2(new_n702_), .ZN(new_n739_));
  AND4_X1   g538(.A1(new_n704_), .A2(new_n739_), .A3(KEYINPUT44), .A4(new_n685_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n704_), .B1(new_n703_), .B2(KEYINPUT44), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n734_), .B(KEYINPUT103), .C1(new_n740_), .C2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G50gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT103), .B1(new_n706_), .B2(new_n734_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n730_), .B1(new_n738_), .B2(new_n746_), .ZN(G1331gat));
  NAND2_X1  g546(.A1(new_n654_), .A2(new_n514_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n748_), .A2(new_n655_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n653_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(G57gat), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n658_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n479_), .A2(new_n513_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT106), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(KEYINPUT106), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NOR4_X1   g555(.A1(new_n756_), .A2(new_n593_), .A3(new_n655_), .A4(new_n696_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n640_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n751_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT107), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n758_), .A2(new_n761_), .A3(new_n751_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n752_), .B1(new_n760_), .B2(new_n762_), .ZN(G1332gat));
  INV_X1    g562(.A(G64gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n757_), .A2(new_n764_), .A3(new_n475_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G64gat), .B1(new_n750_), .B2(new_n456_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT48), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT108), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n765_), .A2(new_n770_), .A3(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1333gat));
  INV_X1    g571(.A(G71gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n757_), .A2(new_n773_), .A3(new_n419_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G71gat), .B1(new_n750_), .B2(new_n478_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(KEYINPUT49), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(KEYINPUT49), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n774_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n774_), .B(KEYINPUT109), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(G1334gat));
  NAND3_X1  g581(.A1(new_n757_), .A2(new_n273_), .A3(new_n673_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G78gat), .B1(new_n750_), .B2(new_n674_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT50), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT110), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n783_), .A2(new_n788_), .A3(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1335gat));
  INV_X1    g589(.A(G85gat), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n748_), .A2(new_n607_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n739_), .A2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT111), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n791_), .B1(new_n794_), .B2(new_n640_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n754_), .A2(new_n755_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n681_), .A2(new_n593_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n798_), .A2(G85gat), .A3(new_n658_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n795_), .A2(new_n799_), .ZN(G1336gat));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n456_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n802_));
  OR3_X1    g601(.A1(new_n801_), .A2(new_n802_), .A3(G92gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(G92gat), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n475_), .A2(G92gat), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n803_), .A2(new_n804_), .B1(new_n794_), .B2(new_n805_), .ZN(G1337gat));
  AOI21_X1  g605(.A(new_n520_), .B1(new_n794_), .B2(new_n419_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n419_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n798_), .A2(new_n808_), .ZN(new_n809_));
  OR3_X1    g608(.A1(new_n807_), .A2(KEYINPUT51), .A3(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT51), .B1(new_n807_), .B2(new_n809_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1338gat));
  XNOR2_X1  g611(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n739_), .A2(new_n792_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n282_), .B1(new_n814_), .B2(new_n474_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT52), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n793_), .A2(new_n289_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n282_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n289_), .A2(G106gat), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n797_), .B(new_n821_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT113), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n813_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n824_));
  AND4_X1   g623(.A1(new_n823_), .A2(new_n819_), .A3(new_n816_), .A4(new_n813_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1339gat));
  NAND4_X1  g625(.A1(new_n497_), .A2(G229gat), .A3(G233gat), .A4(new_n501_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n504_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n509_), .B1(new_n828_), .B2(new_n498_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n506_), .A2(new_n509_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n590_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n580_), .A2(new_n574_), .A3(new_n582_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n588_), .A2(KEYINPUT55), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n589_), .B1(new_n583_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n831_), .B1(KEYINPUT56), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n833_), .A2(new_n835_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT117), .B1(new_n689_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n836_), .A2(KEYINPUT56), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n843_), .A2(new_n590_), .A3(new_n839_), .A4(new_n830_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n696_), .A2(new_n842_), .A3(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n837_), .A2(KEYINPUT58), .A3(new_n839_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n841_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n590_), .A2(new_n513_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n590_), .A2(KEYINPUT115), .A3(new_n513_), .ZN(new_n853_));
  OR2_X1    g652(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n833_), .A2(new_n835_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n852_), .B(new_n853_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n584_), .A2(new_n590_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n830_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(new_n860_), .B2(new_n650_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n862_), .B(new_n680_), .C1(new_n857_), .C2(new_n859_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n607_), .B1(new_n849_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n655_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n514_), .A4(new_n593_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT54), .B1(new_n638_), .B2(new_n513_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n865_), .A2(new_n870_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n373_), .A2(new_n658_), .A3(new_n478_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(KEYINPUT118), .Z(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT59), .ZN(new_n875_));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875_), .B2(new_n514_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n874_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n397_), .A3(new_n513_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1340gat));
  OAI21_X1  g678(.A(G120gat), .B1(new_n875_), .B2(new_n593_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n395_), .B1(new_n593_), .B2(KEYINPUT60), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n877_), .B(new_n881_), .C1(KEYINPUT60), .C2(new_n395_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1341gat));
  OAI21_X1  g682(.A(G127gat), .B1(new_n875_), .B2(new_n655_), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n874_), .A2(G127gat), .A3(new_n655_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1342gat));
  OAI21_X1  g685(.A(G134gat), .B1(new_n875_), .B2(new_n689_), .ZN(new_n887_));
  OR3_X1    g686(.A1(new_n874_), .A2(G134gat), .A3(new_n651_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1343gat));
  NOR4_X1   g688(.A1(new_n658_), .A2(new_n475_), .A3(new_n289_), .A4(new_n419_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n871_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n513_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n654_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g694(.A1(new_n871_), .A2(new_n607_), .A3(new_n890_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT61), .B(G155gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n896_), .B(KEYINPUT119), .ZN(new_n901_));
  INV_X1    g700(.A(new_n899_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(new_n903_), .ZN(G1346gat));
  AOI21_X1  g703(.A(G162gat), .B1(new_n891_), .B2(new_n652_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n689_), .A2(new_n233_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT120), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n891_), .B2(new_n907_), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n456_), .A2(new_n454_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n513_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n674_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n911_), .B2(new_n910_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n315_), .B1(new_n871_), .B2(new_n913_), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT62), .Z(new_n915_));
  NOR3_X1   g714(.A1(new_n673_), .A2(new_n456_), .A3(new_n454_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n871_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(new_n300_), .A3(new_n513_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n915_), .A2(new_n919_), .ZN(G1348gat));
  OAI21_X1  g719(.A(new_n301_), .B1(new_n917_), .B2(new_n593_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n289_), .B1(new_n865_), .B2(new_n870_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  OAI211_X1 g723(.A(KEYINPUT122), .B(new_n289_), .C1(new_n865_), .C2(new_n870_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n593_), .A2(new_n301_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n924_), .A2(new_n909_), .A3(new_n925_), .A4(new_n926_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n921_), .A2(new_n927_), .ZN(G1349gat));
  NAND4_X1  g727(.A1(new_n924_), .A2(new_n607_), .A3(new_n909_), .A4(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n304_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n309_), .A2(new_n311_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n918_), .A2(new_n931_), .A3(new_n607_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n930_), .A2(KEYINPUT123), .A3(new_n932_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n918_), .A2(new_n312_), .A3(new_n652_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n918_), .A2(new_n696_), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n939_), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n940_));
  AOI21_X1  g739(.A(KEYINPUT124), .B1(new_n939_), .B2(G190gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n938_), .B1(new_n940_), .B2(new_n941_), .ZN(G1351gat));
  OR3_X1    g741(.A1(new_n476_), .A2(KEYINPUT125), .A3(new_n419_), .ZN(new_n943_));
  OAI21_X1  g742(.A(KEYINPUT125), .B1(new_n476_), .B2(new_n419_), .ZN(new_n944_));
  AND3_X1   g743(.A1(new_n943_), .A2(new_n475_), .A3(new_n944_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n871_), .A2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n513_), .ZN(new_n947_));
  OAI21_X1  g746(.A(KEYINPUT126), .B1(new_n947_), .B2(new_n206_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n206_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n946_), .A2(new_n950_), .A3(G197gat), .A4(new_n513_), .ZN(new_n951_));
  AND3_X1   g750(.A1(new_n948_), .A2(new_n949_), .A3(new_n951_), .ZN(G1352gat));
  NAND2_X1  g751(.A1(new_n946_), .A2(new_n654_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g753(.A1(new_n946_), .A2(new_n607_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  AND2_X1   g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n955_), .A2(new_n956_), .A3(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n958_), .B1(new_n955_), .B2(new_n956_), .ZN(G1354gat));
  AOI21_X1  g758(.A(G218gat), .B1(new_n946_), .B2(new_n652_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n696_), .A2(G218gat), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(KEYINPUT127), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n960_), .B1(new_n946_), .B2(new_n962_), .ZN(G1355gat));
endmodule


