//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n966_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n990_, new_n991_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n204_));
  INV_X1    g003(.A(G155gat), .ZN(new_n205_));
  INV_X1    g004(.A(G162gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT3), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT2), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n210_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G141gat), .B(G148gat), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n208_), .A2(KEYINPUT1), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT79), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n208_), .A2(new_n219_), .A3(KEYINPUT1), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n207_), .B(new_n209_), .C1(KEYINPUT1), .C2(new_n208_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n216_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT80), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n225_), .B(new_n216_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n215_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT81), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT81), .B1(new_n227_), .B2(new_n228_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT82), .B(KEYINPUT28), .Z(new_n232_));
  NOR3_X1   g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n232_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n224_), .A2(new_n226_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n215_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n235_), .B1(new_n238_), .B2(KEYINPUT29), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n234_), .B1(new_n239_), .B2(new_n229_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n203_), .B1(new_n233_), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n232_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n239_), .A2(new_n229_), .A3(new_n234_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n202_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT84), .B1(new_n246_), .B2(G204gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT84), .ZN(new_n248_));
  INV_X1    g047(.A(G204gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(G197gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(G204gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(KEYINPUT85), .B(KEYINPUT21), .Z(new_n253_));
  OR2_X1    g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G211gat), .B(G218gat), .Z(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(G197gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n251_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(KEYINPUT21), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n255_), .A2(KEYINPUT21), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n252_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT83), .ZN(new_n264_));
  INV_X1    g063(.A(G106gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT83), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n266_), .B(new_n262_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n265_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G228gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(G78gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n269_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n273_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n264_), .A2(new_n267_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G106gat), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n275_), .B1(new_n277_), .B2(new_n268_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n245_), .B1(new_n274_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n273_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(new_n275_), .A3(new_n268_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n244_), .A4(new_n241_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G127gat), .B(G134gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(G113gat), .B(G120gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n238_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n227_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G225gat), .A2(G233gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G1gat), .B(G29gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(G57gat), .B(G85gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n287_), .A2(KEYINPUT4), .A3(new_n289_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT91), .B(KEYINPUT4), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n238_), .A2(new_n286_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n290_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n291_), .B(new_n296_), .C1(new_n297_), .C2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT33), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n287_), .A2(KEYINPUT4), .A3(new_n289_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n227_), .A2(new_n288_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n300_), .B1(new_n305_), .B2(new_n298_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n296_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT93), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n287_), .A2(new_n308_), .A3(new_n289_), .ZN(new_n309_));
  AOI211_X1 g108(.A(new_n286_), .B(new_n215_), .C1(new_n224_), .C2(new_n226_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT93), .B1(new_n305_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n311_), .A3(new_n300_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n302_), .A2(new_n303_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT23), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G183gat), .A3(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(G183gat), .B2(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT89), .ZN(new_n320_));
  INV_X1    g119(.A(G169gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT22), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT22), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G169gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT88), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n322_), .A2(new_n324_), .A3(KEYINPUT88), .ZN(new_n328_));
  INV_X1    g127(.A(G176gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n318_), .B(new_n331_), .C1(G183gat), .C2(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n320_), .A2(new_n330_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n254_), .A2(new_n258_), .B1(new_n260_), .B2(new_n252_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT25), .B(G183gat), .ZN(new_n336_));
  OR2_X1    g135(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n338_));
  NAND2_X1  g137(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n336_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n317_), .A2(KEYINPUT77), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n315_), .A2(new_n317_), .A3(KEYINPUT77), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n321_), .A2(new_n329_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(KEYINPUT24), .A3(new_n333_), .ZN(new_n346_));
  OR3_X1    g145(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .A4(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n334_), .A2(new_n335_), .A3(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n350_), .A2(KEYINPUT20), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT90), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT19), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n318_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT26), .ZN(new_n357_));
  OR2_X1    g156(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(KEYINPUT75), .A2(G190gat), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n337_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n336_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(G183gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n358_), .A2(new_n364_), .A3(new_n359_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n343_), .A2(new_n344_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n368_));
  AOI21_X1  g167(.A(G176gat), .B1(new_n322_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n368_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n333_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n363_), .B1(new_n367_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n262_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n351_), .A2(new_n352_), .A3(new_n355_), .A4(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n374_), .A2(new_n350_), .A3(KEYINPUT20), .A4(new_n355_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT90), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G8gat), .B(G36gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT18), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT86), .B(KEYINPUT20), .C1(new_n373_), .C2(new_n262_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n334_), .A2(new_n349_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n262_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT20), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n325_), .A2(KEYINPUT76), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n388_), .A2(new_n369_), .B1(G169gat), .B2(G176gat), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n389_), .A2(new_n366_), .B1(new_n356_), .B2(new_n362_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n387_), .B1(new_n390_), .B2(new_n335_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(KEYINPUT86), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n354_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n378_), .A2(new_n382_), .A3(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n376_), .A2(KEYINPUT90), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n376_), .A2(KEYINPUT90), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n393_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n382_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n304_), .A2(new_n300_), .A3(new_n299_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n400_), .A2(KEYINPUT33), .A3(new_n291_), .A4(new_n296_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n313_), .A2(new_n394_), .A3(new_n399_), .A4(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n391_), .A2(KEYINPUT86), .B1(new_n262_), .B2(new_n384_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT20), .B1(new_n373_), .B2(new_n262_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n403_), .A2(new_n406_), .A3(KEYINPUT94), .A4(new_n355_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n386_), .A2(new_n392_), .A3(new_n354_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT94), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n374_), .A2(new_n350_), .A3(KEYINPUT20), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(new_n354_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n407_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n382_), .A2(KEYINPUT32), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n403_), .A2(new_n406_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n375_), .A2(new_n377_), .B1(new_n416_), .B2(new_n354_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n413_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n296_), .B1(new_n400_), .B2(new_n291_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n302_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n415_), .B(new_n418_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n402_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n283_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n279_), .A2(new_n282_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n399_), .A2(new_n394_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n417_), .B2(new_n382_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n382_), .B(KEYINPUT95), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n412_), .A2(new_n428_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n425_), .A2(new_n426_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n420_), .A2(new_n419_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n424_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n423_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n435_), .B(G43gat), .Z(new_n436_));
  NAND2_X1  g235(.A1(new_n373_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n436_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n390_), .A2(new_n438_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n437_), .A2(new_n288_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n288_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(G15gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT30), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n445_), .B(KEYINPUT31), .Z(new_n446_));
  OR3_X1    g245(.A1(new_n440_), .A2(new_n441_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n420_), .A2(new_n419_), .A3(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n279_), .A2(new_n450_), .A3(new_n282_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT96), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n430_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n279_), .A2(new_n450_), .A3(new_n282_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n394_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n382_), .B1(new_n378_), .B2(new_n393_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n426_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n427_), .A2(new_n429_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT96), .B1(new_n454_), .B2(new_n459_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n434_), .A2(new_n449_), .B1(new_n453_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462_));
  INV_X1    g261(.A(G1gat), .ZN(new_n463_));
  INV_X1    g262(.A(G8gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT14), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G1gat), .B(G8gat), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G29gat), .B(G36gat), .Z(new_n469_));
  XOR2_X1   g268(.A(G43gat), .B(G50gat), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n466_), .A2(new_n467_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n468_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n468_), .A2(new_n476_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT15), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n475_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n471_), .A2(KEYINPUT15), .A3(new_n474_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT73), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT73), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n480_), .A2(new_n482_), .A3(new_n486_), .A4(new_n483_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n479_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n475_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n480_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n477_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n478_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G113gat), .B(G141gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT74), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G169gat), .B(G197gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n489_), .A2(new_n494_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n494_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n498_), .B1(new_n488_), .B2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n461_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G134gat), .B(G162gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT36), .Z(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT66), .B(KEYINPUT34), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G232gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT35), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT64), .ZN(new_n515_));
  AND2_X1   g314(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT10), .ZN(new_n519_));
  INV_X1    g318(.A(G99gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(KEYINPUT64), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n265_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT6), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(G99gat), .A3(G106gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(G85gat), .ZN(new_n531_));
  INV_X1    g330(.A(G92gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(KEYINPUT9), .A3(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(KEYINPUT9), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n530_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n525_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n533_), .A2(new_n534_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI211_X1 g342(.A(KEYINPUT8), .B(new_n539_), .C1(new_n543_), .C2(new_n530_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT8), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT7), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(new_n520_), .A3(new_n265_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n530_), .A2(new_n540_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n539_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n545_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n538_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(KEYINPUT68), .B(new_n514_), .C1(new_n551_), .C2(new_n490_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n511_), .A2(KEYINPUT35), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT67), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(G106gat), .B1(new_n518_), .B2(new_n523_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n530_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n527_), .A2(new_n529_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n547_), .A2(new_n540_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n549_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT8), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n548_), .A2(new_n545_), .A3(new_n549_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n559_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n565_), .A2(new_n475_), .B1(new_n513_), .B2(new_n512_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT65), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(KEYINPUT65), .A3(new_n564_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n559_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n482_), .A2(new_n483_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n566_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n556_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(new_n569_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n538_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n571_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n555_), .B1(new_n577_), .B2(new_n566_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n508_), .B1(new_n573_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n556_), .A2(new_n572_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(new_n566_), .A3(new_n555_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n507_), .A2(KEYINPUT36), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n580_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n579_), .A2(KEYINPUT37), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT69), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n508_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT69), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n583_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT37), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n585_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT17), .ZN(new_n594_));
  XOR2_X1   g393(.A(G127gat), .B(G155gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT70), .B(KEYINPUT16), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G57gat), .B(G64gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G71gat), .B(G78gat), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(KEYINPUT11), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(KEYINPUT11), .ZN(new_n603_));
  INV_X1    g402(.A(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n600_), .A2(KEYINPUT11), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(G231gat), .ZN(new_n608_));
  INV_X1    g407(.A(G233gat), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n468_), .A2(new_n476_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n468_), .B2(new_n476_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n607_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n614_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n607_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n612_), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n599_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT71), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n599_), .ZN(new_n622_));
  OAI22_X1  g421(.A1(new_n594_), .A2(new_n619_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n615_), .A2(new_n618_), .ZN(new_n624_));
  OAI211_X1 g423(.A(KEYINPUT17), .B(new_n599_), .C1(new_n624_), .C2(new_n620_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n565_), .A2(new_n607_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n607_), .B(new_n538_), .C1(new_n544_), .C2(new_n550_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n628_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT12), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n565_), .B2(new_n607_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n617_), .A2(KEYINPUT12), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n634_), .B(new_n630_), .C1(new_n570_), .C2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n636_), .B2(new_n628_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT5), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n639_), .B(new_n640_), .Z(new_n641_));
  NAND2_X1  g440(.A1(new_n637_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n635_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n575_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT12), .B1(new_n551_), .B2(new_n617_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n631_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n627_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n641_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(new_n632_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n642_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT13), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n642_), .A2(KEYINPUT13), .A3(new_n649_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n593_), .A2(new_n626_), .A3(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT72), .Z(new_n656_));
  NAND4_X1  g455(.A1(new_n504_), .A2(new_n656_), .A3(new_n463_), .A4(new_n431_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT38), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n659_));
  INV_X1    g458(.A(new_n503_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n654_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n626_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT97), .ZN(new_n665_));
  INV_X1    g464(.A(new_n591_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n461_), .B2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n431_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n283_), .A2(new_n422_), .B1(new_n668_), .B2(new_n430_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n449_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n452_), .B1(new_n451_), .B2(new_n430_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n454_), .A2(new_n459_), .A3(KEYINPUT96), .ZN(new_n672_));
  OAI22_X1  g471(.A1(new_n669_), .A2(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(KEYINPUT97), .A3(new_n591_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n664_), .B1(new_n667_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n431_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n659_), .B1(new_n676_), .B2(G1gat), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT98), .B(new_n463_), .C1(new_n675_), .C2(new_n431_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n658_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(G1324gat));
  AND2_X1   g480(.A1(new_n504_), .A2(new_n656_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n464_), .A3(new_n459_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n464_), .B1(new_n675_), .B2(new_n459_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n684_), .A2(new_n685_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT40), .B(new_n683_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1325gat));
  INV_X1    g491(.A(new_n675_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G15gat), .B1(new_n693_), .B2(new_n449_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n695_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n682_), .A2(new_n443_), .A3(new_n670_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n696_), .A2(new_n697_), .A3(new_n698_), .ZN(G1326gat));
  INV_X1    g498(.A(G22gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n682_), .A2(new_n700_), .A3(new_n424_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G22gat), .B1(new_n693_), .B2(new_n283_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(KEYINPUT42), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(KEYINPUT42), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n701_), .B1(new_n703_), .B2(new_n704_), .ZN(G1327gat));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n654_), .A2(new_n662_), .A3(new_n660_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(new_n461_), .B2(new_n593_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n583_), .B1(new_n579_), .B2(new_n586_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n589_), .A2(KEYINPUT69), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n592_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n584_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n673_), .A2(new_n717_), .A3(new_n708_), .ZN(new_n718_));
  AOI211_X1 g517(.A(new_n706_), .B(new_n707_), .C1(new_n713_), .C2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n431_), .A2(G29gat), .ZN(new_n720_));
  INV_X1    g519(.A(new_n707_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n461_), .A2(new_n593_), .A3(new_n709_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n711_), .B1(new_n673_), .B2(new_n717_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(new_n706_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n707_), .B1(new_n713_), .B2(new_n718_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT103), .B1(new_n727_), .B2(KEYINPUT44), .ZN(new_n728_));
  AOI211_X1 g527(.A(new_n719_), .B(new_n720_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n654_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n666_), .A2(new_n662_), .ZN(new_n731_));
  NOR4_X1   g530(.A1(new_n461_), .A2(new_n503_), .A3(new_n730_), .A4(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G29gat), .B1(new_n732_), .B2(new_n431_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT104), .B1(new_n729_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n735_));
  INV_X1    g534(.A(new_n733_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n726_), .A2(new_n728_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n727_), .A2(KEYINPUT44), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n735_), .B(new_n736_), .C1(new_n739_), .C2(new_n720_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n734_), .A2(new_n740_), .ZN(G1328gat));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  INV_X1    g541(.A(G36gat), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n719_), .A2(new_n430_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n737_), .B2(new_n744_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n430_), .A2(KEYINPUT105), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n430_), .A2(KEYINPUT105), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n732_), .A2(new_n743_), .A3(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n742_), .B1(new_n745_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n752_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n738_), .A2(new_n459_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n728_), .B2(new_n726_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT46), .B(new_n754_), .C1(new_n756_), .C2(new_n743_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n753_), .A2(new_n757_), .ZN(G1329gat));
  NAND2_X1  g557(.A1(new_n670_), .A2(G43gat), .ZN(new_n759_));
  AOI211_X1 g558(.A(new_n719_), .B(new_n759_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G43gat), .B1(new_n732_), .B2(new_n670_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT47), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n763_));
  INV_X1    g562(.A(new_n761_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n763_), .B(new_n764_), .C1(new_n739_), .C2(new_n759_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1330gat));
  INV_X1    g565(.A(G50gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n732_), .A2(new_n767_), .A3(new_n424_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n283_), .B1(new_n727_), .B2(KEYINPUT44), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n769_), .B(new_n767_), .C1(new_n737_), .C2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n725_), .B1(new_n724_), .B2(new_n706_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n727_), .A2(KEYINPUT103), .A3(KEYINPUT44), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT107), .B1(new_n774_), .B2(G50gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n768_), .B1(new_n771_), .B2(new_n775_), .ZN(G1331gat));
  NOR2_X1   g575(.A1(new_n461_), .A2(new_n660_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n717_), .A2(new_n662_), .A3(new_n654_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n780_), .A2(KEYINPUT108), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n431_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(KEYINPUT108), .ZN(new_n783_));
  AOI21_X1  g582(.A(G57gat), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n503_), .A2(new_n626_), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n654_), .B(new_n785_), .C1(new_n667_), .C2(new_n674_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(G57gat), .A3(new_n431_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n787_), .A2(KEYINPUT109), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n787_), .A2(KEYINPUT109), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n784_), .A2(new_n788_), .A3(new_n789_), .ZN(G1332gat));
  INV_X1    g589(.A(G64gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n780_), .A2(new_n791_), .A3(new_n749_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT48), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n786_), .A2(new_n749_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(G64gat), .ZN(new_n795_));
  AOI211_X1 g594(.A(KEYINPUT48), .B(new_n791_), .C1(new_n786_), .C2(new_n749_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(G1333gat));
  OR3_X1    g596(.A1(new_n779_), .A2(G71gat), .A3(new_n449_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n786_), .A2(new_n670_), .ZN(new_n799_));
  XOR2_X1   g598(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(G71gat), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n799_), .B2(G71gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(G1334gat));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n786_), .A2(new_n424_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(G78gat), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT50), .B(new_n272_), .C1(new_n786_), .C2(new_n424_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n424_), .A2(new_n272_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT111), .ZN(new_n809_));
  OAI22_X1  g608(.A1(new_n806_), .A2(new_n807_), .B1(new_n779_), .B2(new_n809_), .ZN(G1335gat));
  NOR2_X1   g609(.A1(new_n731_), .A2(new_n654_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n777_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G85gat), .B1(new_n812_), .B2(new_n431_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n654_), .A2(new_n626_), .A3(new_n660_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT112), .B1(new_n722_), .B2(new_n723_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n713_), .A2(new_n718_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n815_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n431_), .A2(G85gat), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT113), .Z(new_n821_));
  AOI21_X1  g620(.A(new_n813_), .B1(new_n819_), .B2(new_n821_), .ZN(G1336gat));
  AOI21_X1  g621(.A(new_n532_), .B1(new_n819_), .B2(new_n749_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n812_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n824_), .A2(G92gat), .A3(new_n430_), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n823_), .A2(KEYINPUT114), .A3(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n823_), .B2(new_n825_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(G1337gat));
  AOI21_X1  g627(.A(new_n520_), .B1(new_n819_), .B2(new_n670_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n812_), .A2(new_n670_), .A3(new_n524_), .ZN(new_n830_));
  OR3_X1    g629(.A1(new_n829_), .A2(KEYINPUT51), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT51), .B1(new_n829_), .B2(new_n830_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1338gat));
  NAND3_X1  g632(.A1(new_n812_), .A2(new_n265_), .A3(new_n424_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n814_), .A2(new_n424_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n713_), .B2(new_n718_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n265_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n836_), .A2(KEYINPUT52), .A3(new_n265_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n834_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g641(.A1(new_n459_), .A2(new_n432_), .A3(new_n449_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n660_), .A2(new_n649_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n636_), .B2(new_n628_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n636_), .A2(new_n628_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n636_), .A2(new_n845_), .A3(new_n628_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n641_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n627_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n647_), .B1(new_n853_), .B2(new_n845_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n849_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(KEYINPUT56), .A3(new_n641_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n844_), .B1(new_n852_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n485_), .A2(new_n487_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(new_n477_), .A3(new_n493_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n499_), .B1(new_n492_), .B2(new_n478_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n500_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n649_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n648_), .B1(new_n647_), .B2(new_n632_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT117), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n650_), .A2(new_n868_), .A3(new_n863_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n591_), .B1(new_n858_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT118), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n873_), .B(new_n591_), .C1(new_n858_), .C2(new_n870_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n872_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n863_), .A2(new_n649_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n852_), .B2(new_n857_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT58), .ZN(new_n879_));
  INV_X1    g678(.A(new_n877_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT56), .B1(new_n856_), .B2(new_n641_), .ZN(new_n881_));
  AOI211_X1 g680(.A(new_n851_), .B(new_n648_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n593_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n844_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n650_), .A2(new_n868_), .A3(new_n863_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n868_), .B1(new_n650_), .B2(new_n863_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n666_), .B1(new_n887_), .B2(new_n890_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n879_), .A2(new_n885_), .B1(new_n891_), .B2(KEYINPUT57), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n626_), .B1(new_n876_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n785_), .A2(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n503_), .A2(KEYINPUT115), .A3(new_n626_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n654_), .A2(new_n894_), .A3(new_n896_), .A4(new_n897_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n896_), .A2(new_n653_), .A3(new_n652_), .A4(new_n897_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT116), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n717_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT54), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n283_), .B(new_n843_), .C1(new_n893_), .C2(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT59), .ZN(new_n904_));
  INV_X1    g703(.A(G113gat), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n904_), .A2(new_n905_), .A3(new_n503_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(KEYINPUT120), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n901_), .B(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT57), .B(new_n591_), .C1(new_n858_), .C2(new_n870_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n717_), .B1(new_n878_), .B2(KEYINPUT58), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n883_), .A2(new_n884_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n875_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n871_), .B2(KEYINPUT118), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n874_), .B2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n909_), .B1(new_n916_), .B2(new_n626_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n917_), .A2(new_n918_), .A3(new_n283_), .A4(new_n843_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n907_), .A2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n905_), .B1(new_n920_), .B2(new_n503_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  OAI211_X1 g722(.A(KEYINPUT121), .B(new_n905_), .C1(new_n920_), .C2(new_n503_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n906_), .B1(new_n923_), .B2(new_n924_), .ZN(G1340gat));
  OAI21_X1  g724(.A(G120gat), .B1(new_n904_), .B2(new_n654_), .ZN(new_n926_));
  INV_X1    g725(.A(G120gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n654_), .B2(KEYINPUT60), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(KEYINPUT60), .B2(new_n927_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n926_), .B1(new_n920_), .B2(new_n929_), .ZN(G1341gat));
  OR3_X1    g729(.A1(new_n920_), .A2(G127gat), .A3(new_n662_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G127gat), .B1(new_n904_), .B2(new_n662_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1342gat));
  OR3_X1    g732(.A1(new_n920_), .A2(G134gat), .A3(new_n591_), .ZN(new_n934_));
  OAI21_X1  g733(.A(G134gat), .B1(new_n904_), .B2(new_n593_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1343gat));
  AND2_X1   g735(.A1(new_n917_), .A2(new_n449_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n749_), .A2(new_n432_), .A3(new_n283_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n937_), .A2(new_n660_), .A3(new_n938_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g739(.A1(new_n937_), .A2(new_n938_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n654_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT122), .B(G148gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1345gat));
  NOR2_X1   g743(.A1(new_n941_), .A2(new_n662_), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT61), .B(G155gat), .Z(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(G1346gat));
  OAI21_X1  g746(.A(G162gat), .B1(new_n941_), .B2(new_n593_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n666_), .A2(new_n206_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n941_), .B2(new_n949_), .ZN(G1347gat));
  NOR3_X1   g749(.A1(new_n748_), .A2(new_n431_), .A3(new_n449_), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n283_), .B(new_n951_), .C1(new_n893_), .C2(new_n902_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n953_), .A2(new_n327_), .A3(new_n328_), .A4(new_n660_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n951_), .A2(new_n660_), .ZN(new_n956_));
  XOR2_X1   g755(.A(new_n956_), .B(KEYINPUT123), .Z(new_n957_));
  AND2_X1   g756(.A1(new_n917_), .A2(new_n283_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n955_), .B1(new_n959_), .B2(G169gat), .ZN(new_n960_));
  AOI211_X1 g759(.A(KEYINPUT62), .B(new_n321_), .C1(new_n957_), .C2(new_n958_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n954_), .B1(new_n960_), .B2(new_n961_), .ZN(G1348gat));
  NOR2_X1   g761(.A1(new_n952_), .A2(new_n654_), .ZN(new_n963_));
  XOR2_X1   g762(.A(KEYINPUT124), .B(G176gat), .Z(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1349gat));
  NOR2_X1   g764(.A1(new_n952_), .A2(new_n662_), .ZN(new_n966_));
  MUX2_X1   g765(.A(G183gat), .B(new_n336_), .S(new_n966_), .Z(G1350gat));
  OAI211_X1 g766(.A(new_n953_), .B(new_n666_), .C1(new_n341_), .C2(new_n340_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969_));
  OAI211_X1 g768(.A(new_n969_), .B(G190gat), .C1(new_n952_), .C2(new_n593_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  NAND4_X1  g770(.A1(new_n917_), .A2(new_n283_), .A3(new_n717_), .A4(new_n951_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n969_), .B1(new_n972_), .B2(G190gat), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n968_), .B1(new_n971_), .B2(new_n973_), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n974_), .A2(new_n975_), .ZN(new_n976_));
  OAI211_X1 g775(.A(KEYINPUT126), .B(new_n968_), .C1(new_n971_), .C2(new_n973_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(G1351gat));
  NOR3_X1   g777(.A1(new_n748_), .A2(new_n431_), .A3(new_n283_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n937_), .A2(new_n979_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n980_), .A2(new_n503_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(new_n246_), .ZN(G1352gat));
  NOR2_X1   g781(.A1(new_n980_), .A2(new_n654_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(new_n983_), .B(new_n249_), .ZN(G1353gat));
  NOR2_X1   g783(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n985_), .B1(new_n980_), .B2(new_n662_), .ZN(new_n986_));
  XOR2_X1   g785(.A(KEYINPUT63), .B(G211gat), .Z(new_n987_));
  NAND4_X1  g786(.A1(new_n937_), .A2(new_n626_), .A3(new_n979_), .A4(new_n987_), .ZN(new_n988_));
  AND2_X1   g787(.A1(new_n986_), .A2(new_n988_), .ZN(G1354gat));
  OAI21_X1  g788(.A(G218gat), .B1(new_n980_), .B2(new_n593_), .ZN(new_n990_));
  OR2_X1    g789(.A1(new_n591_), .A2(G218gat), .ZN(new_n991_));
  OAI21_X1  g790(.A(new_n990_), .B1(new_n980_), .B2(new_n991_), .ZN(G1355gat));
endmodule


