//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203_));
  INV_X1    g002(.A(G78gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G71gat), .ZN(new_n205_));
  INV_X1    g004(.A(G71gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G78gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209_));
  INV_X1    g008(.A(G57gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(G64gat), .ZN(new_n211_));
  INV_X1    g010(.A(G64gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(G57gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n209_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(G57gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(G64gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT68), .ZN(new_n217_));
  AOI211_X1 g016(.A(new_n203_), .B(new_n208_), .C1(new_n214_), .C2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n208_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n217_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(KEYINPUT11), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n214_), .A2(new_n203_), .A3(new_n217_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n218_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT67), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(KEYINPUT6), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT6), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT66), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n228_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT7), .ZN(new_n234_));
  INV_X1    g033(.A(G99gat), .ZN(new_n235_));
  INV_X1    g034(.A(G106gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n224_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n231_), .A2(KEYINPUT66), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n229_), .A2(KEYINPUT6), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(G99gat), .A4(G106gat), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n227_), .A2(new_n233_), .A3(new_n239_), .A4(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G85gat), .B(G92gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT8), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n228_), .A2(new_n231_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n237_), .A2(new_n248_), .A3(new_n224_), .A4(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n244_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT8), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n248_), .A2(new_n249_), .ZN(new_n254_));
  OR2_X1    g053(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n255_));
  OR2_X1    g054(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(G85gat), .B(G92gat), .C1(KEYINPUT65), .C2(KEYINPUT9), .ZN(new_n260_));
  OAI211_X1 g059(.A(KEYINPUT65), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n260_), .A2(new_n261_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n254_), .B(new_n259_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n247_), .A2(new_n253_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n223_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n223_), .A2(new_n265_), .A3(KEYINPUT70), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n223_), .B2(new_n265_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n217_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT68), .B1(new_n215_), .B2(new_n216_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT11), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(new_n222_), .A3(new_n208_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n220_), .A2(KEYINPUT11), .A3(new_n219_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n253_), .A2(new_n264_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n277_), .A2(new_n279_), .A3(KEYINPUT69), .A4(new_n247_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n268_), .A2(new_n269_), .A3(new_n271_), .A4(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G230gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n266_), .A2(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n233_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n245_), .B1(new_n287_), .B2(new_n227_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(new_n278_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n283_), .B1(new_n289_), .B2(new_n277_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n223_), .A2(new_n265_), .A3(KEYINPUT12), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G120gat), .B(G148gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(G176gat), .B(G204gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n284_), .A2(new_n292_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n297_), .B1(new_n284_), .B2(new_n292_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI211_X1 g101(.A(new_n299_), .B(new_n297_), .C1(new_n284_), .C2(new_n292_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n202_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n301_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(new_n299_), .A3(new_n298_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n303_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT13), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G29gat), .B(G36gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G43gat), .B(G50gat), .Z(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G43gat), .B(G50gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT76), .B(G15gat), .ZN(new_n318_));
  INV_X1    g117(.A(G22gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G1gat), .B(G8gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G1gat), .A2(G8gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT14), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n320_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n323_), .B1(new_n325_), .B2(new_n320_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n317_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n320_), .A2(new_n325_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n323_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n314_), .A2(new_n316_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT15), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT15), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n317_), .A2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n332_), .A2(new_n334_), .A3(new_n326_), .A4(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G229gat), .A2(G233gat), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n329_), .A2(new_n337_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n329_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT79), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n332_), .A2(new_n326_), .A3(new_n333_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n339_), .B1(new_n329_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n340_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G113gat), .B(G141gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT81), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT82), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G169gat), .B(G197gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT80), .B1(new_n350_), .B2(KEYINPUT83), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n345_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n345_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n352_), .B1(new_n355_), .B2(new_n350_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT19), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT97), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT21), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G197gat), .B(G204gat), .Z(new_n364_));
  OR2_X1    g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n363_), .B(new_n364_), .C1(KEYINPUT21), .C2(new_n361_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n369_));
  INV_X1    g168(.A(G183gat), .ZN(new_n370_));
  INV_X1    g169(.A(G190gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT23), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(G183gat), .A3(G190gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n369_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT86), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(G183gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT84), .ZN(new_n381_));
  OR3_X1    g180(.A1(new_n370_), .A2(KEYINPUT85), .A3(KEYINPUT25), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT26), .B(G190gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT85), .B1(new_n370_), .B2(KEYINPUT25), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  OAI221_X1 g184(.A(new_n375_), .B1(new_n377_), .B2(new_n378_), .C1(new_n381_), .C2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT22), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT87), .B1(new_n387_), .B2(G169gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(G176gat), .B1(new_n387_), .B2(G169gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n390_));
  INV_X1    g189(.A(G169gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(KEYINPUT22), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n377_), .B1(new_n393_), .B2(KEYINPUT88), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n372_), .A2(KEYINPUT89), .A3(new_n374_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n396_), .B(KEYINPUT23), .C1(new_n370_), .C2(new_n371_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n395_), .B(new_n397_), .C1(G183gat), .C2(G190gat), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n394_), .B(new_n398_), .C1(KEYINPUT88), .C2(new_n393_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n368_), .A2(new_n386_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT20), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n372_), .A2(new_n374_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(G183gat), .B2(G190gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT100), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n377_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT86), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n376_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT100), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT22), .B(G169gat), .ZN(new_n409_));
  INV_X1    g208(.A(G176gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n403_), .A2(new_n405_), .A3(new_n408_), .A4(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n378_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n369_), .B1(new_n413_), .B2(new_n376_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT25), .B(G183gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n383_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n414_), .A2(new_n416_), .A3(new_n395_), .A4(new_n397_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n401_), .B1(new_n418_), .B2(new_n367_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n360_), .B1(new_n400_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT101), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT104), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT18), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n425_), .B(new_n426_), .Z(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT20), .B1(new_n418_), .B2(new_n367_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(new_n359_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n399_), .A2(new_n386_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n367_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n422_), .A2(new_n423_), .A3(new_n427_), .A4(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n427_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n428_), .A2(KEYINPUT102), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT102), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n436_), .B(KEYINPUT20), .C1(new_n418_), .C2(new_n367_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n431_), .A3(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n438_), .A2(KEYINPUT103), .A3(new_n359_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n400_), .A2(new_n419_), .A3(new_n360_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n438_), .A2(new_n359_), .B1(KEYINPUT103), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n434_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n420_), .A2(new_n421_), .ZN(new_n443_));
  AOI211_X1 g242(.A(KEYINPUT101), .B(new_n360_), .C1(new_n400_), .C2(new_n419_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n427_), .B(new_n432_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT104), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n433_), .A2(new_n442_), .A3(new_n446_), .A4(KEYINPUT27), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n432_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n434_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n445_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT27), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G127gat), .B(G134gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G113gat), .B(G120gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G155gat), .A2(G162gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT96), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G141gat), .A2(G148gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT3), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n462_), .A2(new_n463_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n461_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT1), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT95), .B1(new_n459_), .B2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n460_), .B1(new_n459_), .B2(new_n472_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT95), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n458_), .A2(new_n475_), .A3(KEYINPUT1), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n473_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n465_), .B(KEYINPUT94), .Z(new_n478_));
  INV_X1    g277(.A(KEYINPUT2), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n477_), .A2(new_n478_), .B1(new_n479_), .B2(new_n461_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT93), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n471_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n457_), .A2(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n471_), .B(new_n455_), .C1(new_n480_), .C2(new_n482_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(KEYINPUT4), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G225gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT4), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n457_), .A2(new_n489_), .A3(new_n483_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G1gat), .B(G29gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(G85gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT0), .B(G57gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n491_), .A2(new_n492_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n447_), .A2(new_n452_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G227gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(new_n206_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G15gat), .B(G43gat), .Z(new_n506_));
  NAND3_X1  g305(.A1(new_n399_), .A2(KEYINPUT30), .A3(new_n386_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT30), .B1(new_n399_), .B2(new_n386_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n430_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n506_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n507_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n510_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n511_), .B1(new_n510_), .B2(new_n515_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n505_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n518_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n505_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n457_), .B(KEYINPUT31), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G99gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n519_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n480_), .A2(new_n482_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT29), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .A4(new_n471_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT28), .B1(new_n483_), .B2(KEYINPUT29), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G22gat), .B(G50gat), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n368_), .B1(new_n483_), .B2(KEYINPUT29), .ZN(new_n538_));
  OAI211_X1 g337(.A(G228gat), .B(G233gat), .C1(new_n368_), .C2(KEYINPUT98), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(KEYINPUT99), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G78gat), .B(G106gat), .Z(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n538_), .B(new_n539_), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n532_), .A2(new_n533_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n534_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n542_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n544_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n541_), .A2(new_n543_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n541_), .B1(new_n543_), .B2(new_n551_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n527_), .B(new_n528_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT99), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n537_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n550_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n541_), .A2(new_n543_), .A3(new_n551_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n519_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n525_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n559_), .B(new_n560_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n503_), .B1(new_n554_), .B2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n552_), .A2(new_n553_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n427_), .A2(KEYINPUT32), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n422_), .A2(new_n432_), .A3(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n439_), .A2(new_n441_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n501_), .B(new_n567_), .C1(new_n568_), .C2(new_n566_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n486_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n484_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n497_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT33), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n500_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n491_), .A2(KEYINPUT33), .A3(new_n492_), .A4(new_n499_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n574_), .A2(new_n445_), .A3(new_n449_), .A4(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n569_), .A2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n561_), .A2(new_n562_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n565_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n357_), .B1(new_n564_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT105), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n310_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n564_), .A2(new_n579_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(KEYINPUT105), .A3(new_n357_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G190gat), .B(G218gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT74), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n589_), .A2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n594_), .A2(KEYINPUT35), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(KEYINPUT35), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n289_), .A2(new_n333_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n334_), .A2(new_n336_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n265_), .ZN(new_n599_));
  AOI211_X1 g398(.A(new_n595_), .B(new_n596_), .C1(new_n597_), .C2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT75), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n597_), .A2(new_n599_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n595_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n600_), .A2(KEYINPUT75), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n591_), .B(new_n592_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n600_), .A2(KEYINPUT75), .B1(new_n603_), .B2(new_n595_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n590_), .A4(new_n589_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n607_), .A2(KEYINPUT37), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT37), .B1(new_n607_), .B2(new_n610_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n223_), .B(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n327_), .A2(new_n328_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n277_), .B(new_n614_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT78), .ZN(new_n622_));
  XOR2_X1   g421(.A(G127gat), .B(G155gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT16), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT17), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n621_), .A2(new_n622_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT17), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n618_), .A2(new_n620_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n622_), .B1(new_n621_), .B2(new_n627_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n613_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n585_), .A2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n637_), .A2(G1gat), .A3(new_n502_), .ZN(new_n638_));
  XOR2_X1   g437(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n564_), .A2(new_n579_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n607_), .A2(new_n610_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n310_), .A2(new_n635_), .A3(new_n356_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n646_), .B2(new_n502_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n638_), .A2(new_n639_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n640_), .A2(new_n647_), .A3(new_n648_), .ZN(G1324gat));
  NAND2_X1  g448(.A1(new_n447_), .A2(new_n452_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n583_), .A2(new_n642_), .A3(new_n650_), .A4(new_n645_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT107), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT107), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n644_), .A2(new_n653_), .A3(new_n650_), .A4(new_n645_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(G8gat), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT108), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(KEYINPUT39), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n582_), .A2(new_n584_), .A3(new_n636_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n650_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(G8gat), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n655_), .A2(new_n657_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT108), .B(KEYINPUT39), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n652_), .A2(new_n654_), .A3(G8gat), .A4(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(KEYINPUT109), .B(KEYINPUT40), .Z(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT110), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n661_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  OAI21_X1  g467(.A(G15gat), .B1(new_n646_), .B2(new_n578_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT41), .Z(new_n670_));
  OR2_X1    g469(.A1(new_n578_), .A2(G15gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n637_), .B2(new_n671_), .ZN(G1326gat));
  OAI21_X1  g471(.A(G22gat), .B1(new_n646_), .B2(new_n565_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT42), .ZN(new_n674_));
  INV_X1    g473(.A(new_n565_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n658_), .A2(new_n319_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1327gat));
  NOR2_X1   g476(.A1(new_n642_), .A2(new_n634_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n585_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(G29gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n501_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n613_), .B1(new_n564_), .B2(new_n579_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT43), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n684_), .B(new_n613_), .C1(new_n564_), .C2(new_n579_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n309_), .A2(new_n635_), .A3(new_n357_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT44), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n690_), .B(new_n687_), .C1(new_n683_), .C2(new_n685_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT111), .B(new_n680_), .C1(new_n692_), .C2(new_n501_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n694_));
  INV_X1    g493(.A(new_n689_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n691_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n501_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n694_), .B1(new_n697_), .B2(G29gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n681_), .B1(new_n693_), .B2(new_n698_), .ZN(G1328gat));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n692_), .B2(new_n650_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n659_), .A2(G36gat), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n582_), .A2(new_n584_), .A3(new_n678_), .A4(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n700_), .B1(new_n702_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n704_), .B(KEYINPUT45), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n689_), .A2(new_n691_), .A3(new_n659_), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n708_), .B(KEYINPUT46), .C1(new_n701_), .C2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1329gat));
  INV_X1    g510(.A(G43gat), .ZN(new_n712_));
  NOR4_X1   g511(.A1(new_n689_), .A2(new_n691_), .A3(new_n712_), .A4(new_n578_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n578_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n585_), .A2(new_n714_), .A3(new_n678_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(new_n712_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT47), .B1(new_n713_), .B2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n692_), .A2(G43gat), .A3(new_n714_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(new_n712_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n717_), .A2(new_n721_), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n692_), .B2(new_n675_), .ZN(new_n724_));
  AND4_X1   g523(.A1(new_n723_), .A2(new_n585_), .A3(new_n675_), .A4(new_n678_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT112), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n679_), .A2(new_n723_), .A3(new_n675_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n689_), .A2(new_n691_), .A3(new_n565_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n727_), .B(new_n728_), .C1(new_n729_), .C2(new_n723_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n726_), .A2(new_n730_), .ZN(G1331gat));
  NOR3_X1   g530(.A1(new_n641_), .A2(new_n357_), .A3(new_n309_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n636_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(KEYINPUT113), .A3(new_n636_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n210_), .A3(new_n501_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n634_), .A2(new_n356_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n309_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n583_), .A2(new_n642_), .A3(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G57gat), .B1(new_n741_), .B2(new_n502_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(G1332gat));
  NAND4_X1  g542(.A1(new_n735_), .A2(new_n212_), .A3(new_n650_), .A4(new_n736_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G64gat), .B1(new_n741_), .B2(new_n659_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(KEYINPUT48), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n747_), .B(G64gat), .C1(new_n741_), .C2(new_n659_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n744_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT114), .ZN(G1333gat));
  NAND3_X1  g550(.A1(new_n737_), .A2(new_n206_), .A3(new_n714_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G71gat), .B1(new_n741_), .B2(new_n578_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT49), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1334gat));
  NAND3_X1  g554(.A1(new_n737_), .A2(new_n204_), .A3(new_n675_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G78gat), .B1(new_n741_), .B2(new_n565_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT50), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1335gat));
  INV_X1    g558(.A(G85gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n732_), .A2(new_n678_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n502_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT115), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n310_), .A2(new_n635_), .A3(new_n356_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n502_), .A2(new_n760_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n763_), .B1(new_n765_), .B2(new_n766_), .ZN(G1336gat));
  INV_X1    g566(.A(new_n761_), .ZN(new_n768_));
  INV_X1    g567(.A(G92gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n650_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n765_), .A2(new_n650_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n769_), .ZN(G1337gat));
  NAND4_X1  g571(.A1(new_n768_), .A2(new_n255_), .A3(new_n257_), .A4(new_n714_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n765_), .A2(new_n714_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n235_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g575(.A1(new_n768_), .A2(new_n256_), .A3(new_n258_), .A4(new_n675_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n765_), .A2(new_n675_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G106gat), .ZN(new_n780_));
  AOI211_X1 g579(.A(KEYINPUT52), .B(new_n236_), .C1(new_n765_), .C2(new_n675_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n777_), .B(new_n783_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(new_n297_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n289_), .A2(new_n277_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n286_), .A2(new_n291_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n292_), .A2(KEYINPUT55), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n286_), .A2(new_n290_), .A3(new_n793_), .A4(new_n291_), .ZN(new_n794_));
  AOI221_X4 g593(.A(new_n789_), .B1(new_n283_), .B2(new_n791_), .C1(new_n792_), .C2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n794_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n283_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT119), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n788_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n297_), .A2(new_n800_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT120), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n223_), .A2(new_n265_), .A3(KEYINPUT12), .ZN(new_n806_));
  INV_X1    g605(.A(new_n285_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n223_), .B2(new_n265_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n793_), .B1(new_n809_), .B2(new_n290_), .ZN(new_n810_));
  AND4_X1   g609(.A1(new_n793_), .A2(new_n286_), .A3(new_n290_), .A4(new_n291_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n797_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n789_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n796_), .A2(KEYINPUT119), .A3(new_n797_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(KEYINPUT120), .A3(new_n802_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n801_), .A2(new_n805_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n357_), .A2(new_n298_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n329_), .A2(new_n337_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(G229gat), .A3(G233gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n329_), .A2(new_n339_), .A3(new_n343_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n350_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n350_), .B2(new_n345_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n306_), .A2(new_n307_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT57), .B1(new_n827_), .B2(new_n642_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n826_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n642_), .A2(KEYINPUT57), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n825_), .A2(new_n298_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n815_), .B2(new_n788_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n802_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT58), .B(new_n833_), .C1(new_n834_), .C2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n613_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n801_), .A2(new_n803_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n839_), .B2(new_n833_), .ZN(new_n840_));
  OAI22_X1  g639(.A1(new_n830_), .A2(new_n831_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n635_), .B1(new_n828_), .B2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(KEYINPUT118), .A2(KEYINPUT54), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n611_), .A2(new_n612_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n739_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(KEYINPUT117), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847_));
  AOI211_X1 g646(.A(new_n847_), .B(new_n739_), .C1(new_n304_), .C2(new_n308_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n843_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n739_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n302_), .A2(new_n202_), .A3(new_n303_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT13), .B1(new_n306_), .B2(new_n307_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n847_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n845_), .A2(KEYINPUT117), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n856_));
  NAND4_X1  g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n844_), .A4(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n849_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n842_), .A2(new_n858_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n563_), .A2(new_n650_), .A3(new_n502_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(G113gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n357_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n861_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n859_), .A2(KEYINPUT59), .A3(new_n860_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n356_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n868_), .B2(new_n863_), .ZN(G1340gat));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n870_));
  AOI21_X1  g669(.A(G120gat), .B1(new_n310_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT121), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n870_), .B2(G120gat), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n862_), .B(new_n872_), .C1(new_n871_), .C2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n309_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n876_));
  INV_X1    g675(.A(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(G1341gat));
  INV_X1    g677(.A(G127gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n862_), .A2(new_n879_), .A3(new_n634_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n635_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n879_), .ZN(G1342gat));
  INV_X1    g681(.A(G134gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n862_), .A2(new_n883_), .A3(new_n643_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n844_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n883_), .ZN(G1343gat));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n554_), .A2(new_n650_), .A3(new_n502_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n859_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n888_), .ZN(new_n890_));
  AOI211_X1 g689(.A(KEYINPUT122), .B(new_n890_), .C1(new_n842_), .C2(new_n858_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n357_), .B1(new_n889_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G141gat), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n849_), .A2(new_n857_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n830_), .B2(new_n643_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n831_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n804_), .A2(new_n803_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n818_), .B1(new_n898_), .B2(new_n816_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n899_), .B2(new_n829_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n839_), .A2(new_n833_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT58), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n832_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n844_), .B1(new_n904_), .B2(KEYINPUT58), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n896_), .A2(new_n900_), .A3(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n894_), .B1(new_n907_), .B2(new_n635_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT122), .B1(new_n908_), .B2(new_n890_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n827_), .A2(new_n897_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n634_), .B1(new_n910_), .B2(new_n896_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n888_), .B(new_n887_), .C1(new_n911_), .C2(new_n894_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(G141gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n914_), .A3(new_n357_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n893_), .A2(new_n915_), .ZN(G1344gat));
  XNOR2_X1  g715(.A(KEYINPUT123), .B(G148gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n913_), .B2(new_n310_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n917_), .ZN(new_n919_));
  AOI211_X1 g718(.A(new_n309_), .B(new_n919_), .C1(new_n909_), .C2(new_n912_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1345gat));
  OAI21_X1  g720(.A(new_n634_), .B1(new_n889_), .B2(new_n891_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT61), .B(G155gat), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n923_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n913_), .A2(new_n634_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1346gat));
  INV_X1    g726(.A(G162gat), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n913_), .A2(new_n928_), .A3(new_n643_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n844_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n928_), .B2(new_n930_), .ZN(G1347gat));
  XNOR2_X1  g730(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n659_), .A2(new_n563_), .A3(new_n501_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n859_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n356_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n932_), .B1(new_n935_), .B2(new_n391_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n932_), .ZN(new_n937_));
  OAI211_X1 g736(.A(G169gat), .B(new_n937_), .C1(new_n934_), .C2(new_n356_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n935_), .A2(new_n409_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n936_), .A2(new_n938_), .A3(new_n939_), .ZN(G1348gat));
  NOR2_X1   g739(.A1(new_n934_), .A2(new_n309_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(new_n410_), .ZN(G1349gat));
  NOR3_X1   g741(.A1(new_n934_), .A2(new_n635_), .A3(new_n415_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n934_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n634_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n943_), .B1(new_n370_), .B2(new_n945_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n934_), .B2(new_n844_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n643_), .A2(new_n383_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n934_), .B2(new_n948_), .ZN(G1351gat));
  NOR3_X1   g748(.A1(new_n659_), .A2(new_n554_), .A3(new_n501_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n859_), .A2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n951_), .A2(new_n356_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(KEYINPUT125), .B(G197gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n952_), .B(new_n953_), .ZN(G1352gat));
  NOR2_X1   g753(.A1(new_n951_), .A2(new_n309_), .ZN(new_n955_));
  INV_X1    g754(.A(G204gat), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n955_), .B(new_n956_), .ZN(G1353gat));
  INV_X1    g756(.A(new_n951_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n634_), .A2(new_n959_), .ZN(new_n960_));
  XOR2_X1   g759(.A(new_n960_), .B(KEYINPUT126), .Z(new_n961_));
  NOR2_X1   g760(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n961_), .B1(KEYINPUT127), .B2(new_n962_), .ZN(new_n963_));
  OAI211_X1 g762(.A(new_n958_), .B(new_n963_), .C1(KEYINPUT127), .C2(new_n962_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n965_));
  OAI221_X1 g764(.A(new_n965_), .B1(KEYINPUT63), .B2(G211gat), .C1(new_n951_), .C2(new_n961_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n964_), .A2(new_n966_), .ZN(G1354gat));
  OR3_X1    g766(.A1(new_n951_), .A2(G218gat), .A3(new_n642_), .ZN(new_n968_));
  OAI21_X1  g767(.A(G218gat), .B1(new_n951_), .B2(new_n844_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1355gat));
endmodule


