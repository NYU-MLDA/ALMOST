//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n208_));
  OR2_X1    g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(KEYINPUT82), .A3(new_n209_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n203_), .B(new_n206_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(new_n207_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT84), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n203_), .B(KEYINPUT2), .Z(new_n219_));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT83), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n206_), .B(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n218_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n216_), .A2(new_n223_), .A3(KEYINPUT85), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT85), .B1(new_n216_), .B2(new_n223_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT29), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT87), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT88), .B(G197gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(KEYINPUT21), .B(new_n229_), .C1(new_n230_), .C2(G204gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(G211gat), .B(G218gat), .Z(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G204gat), .ZN(new_n234_));
  OR3_X1    g033(.A1(new_n230_), .A2(KEYINPUT90), .A3(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT90), .B1(new_n230_), .B2(new_n234_), .ZN(new_n236_));
  INV_X1    g035(.A(G197gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(G204gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT89), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n231_), .B(new_n233_), .C1(new_n240_), .C2(KEYINPUT21), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(KEYINPUT21), .A3(new_n232_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT91), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(KEYINPUT91), .A3(new_n242_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G228gat), .A2(G233gat), .ZN(new_n248_));
  OAI211_X1 g047(.A(KEYINPUT87), .B(KEYINPUT29), .C1(new_n224_), .C2(new_n225_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n228_), .A2(new_n247_), .A3(new_n248_), .A4(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT92), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n243_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n216_), .A2(new_n223_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT29), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n241_), .A2(KEYINPUT92), .A3(new_n242_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(G228gat), .A3(G233gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(G78gat), .B(G106gat), .Z(new_n258_));
  NAND3_X1  g057(.A1(new_n250_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT85), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n253_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n216_), .A2(new_n223_), .A3(KEYINPUT85), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .A4(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G22gat), .B(G50gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n267_), .A2(new_n271_), .A3(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(KEYINPUT93), .A3(new_n274_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n258_), .B1(new_n250_), .B2(new_n257_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n260_), .A2(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n276_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n277_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n259_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT94), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n278_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n278_), .B2(new_n281_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT18), .B(G64gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(G92gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G8gat), .B(G36gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n291_), .B(KEYINPUT79), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(new_n293_), .ZN(new_n296_));
  INV_X1    g095(.A(G169gat), .ZN(new_n297_));
  INV_X1    g096(.A(G176gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT24), .B1(new_n297_), .B2(new_n298_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n296_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT25), .B(G183gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT26), .B(G190gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n299_), .A2(KEYINPUT24), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n297_), .A2(new_n298_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT22), .B(G169gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(new_n298_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT80), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n292_), .A2(KEYINPUT23), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n295_), .B2(KEYINPUT23), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(G183gat), .B2(G190gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n307_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n246_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT91), .B1(new_n241_), .B2(new_n242_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT19), .ZN(new_n321_));
  INV_X1    g120(.A(new_n243_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT95), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n304_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n303_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT96), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n300_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n299_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n325_), .A2(new_n306_), .A3(new_n328_), .A4(new_n313_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n310_), .B1(new_n296_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n321_), .B1(new_n322_), .B2(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n319_), .A2(KEYINPUT20), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n321_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n245_), .A2(new_n246_), .A3(new_n307_), .A4(new_n315_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT20), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n243_), .B2(new_n332_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n290_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n339_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n321_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n319_), .A2(KEYINPUT20), .A3(new_n334_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n289_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT27), .B1(new_n341_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n344_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n337_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n252_), .A2(new_n255_), .ZN(new_n350_));
  OAI211_X1 g149(.A(KEYINPUT20), .B(new_n319_), .C1(new_n350_), .C2(new_n332_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n349_), .B1(new_n321_), .B2(new_n351_), .ZN(new_n352_));
  MUX2_X1   g151(.A(new_n347_), .B(new_n352_), .S(new_n290_), .Z(new_n353_));
  AOI21_X1  g152(.A(new_n346_), .B1(new_n353_), .B2(KEYINPUT27), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n355_), .B(KEYINPUT98), .Z(new_n356_));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357_));
  INV_X1    g156(.A(G113gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G120gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n262_), .A2(new_n264_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT97), .B1(new_n253_), .B2(new_n360_), .ZN(new_n365_));
  INV_X1    g164(.A(G120gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n359_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT97), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n216_), .A4(new_n223_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n364_), .A2(new_n360_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n356_), .B(new_n363_), .C1(new_n370_), .C2(new_n362_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n356_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT99), .B(KEYINPUT0), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT100), .ZN(new_n375_));
  XOR2_X1   g174(.A(G1gat), .B(G29gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n373_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n316_), .B(new_n360_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G71gat), .B(G99gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT31), .ZN(new_n389_));
  XOR2_X1   g188(.A(G15gat), .B(G43gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G227gat), .A2(G233gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n387_), .B(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n384_), .A2(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n285_), .A2(new_n354_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT101), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n373_), .A2(KEYINPUT33), .A3(new_n380_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n341_), .A3(new_n345_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n356_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n365_), .A2(new_n369_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n362_), .B1(new_n401_), .B2(new_n361_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT4), .B1(new_n364_), .B2(new_n360_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n400_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n370_), .A2(new_n356_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n379_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n382_), .B1(KEYINPUT33), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n397_), .B1(new_n399_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(KEYINPUT33), .ZN(new_n409_));
  INV_X1    g208(.A(new_n382_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n341_), .A2(new_n345_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n411_), .A2(KEYINPUT101), .A3(new_n413_), .A4(new_n398_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n289_), .A2(KEYINPUT32), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n343_), .A2(new_n344_), .A3(new_n415_), .ZN(new_n416_));
  OAI221_X1 g215(.A(new_n416_), .B1(new_n352_), .B2(new_n415_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n408_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n285_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n354_), .B(new_n383_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n396_), .B1(new_n421_), .B2(new_n394_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G232gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT34), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT15), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G43gat), .B(G50gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT73), .B(G29gat), .ZN(new_n430_));
  INV_X1    g229(.A(G36gat), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n431_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n429_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n430_), .A2(new_n431_), .ZN(new_n435_));
  INV_X1    g234(.A(G29gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT73), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT73), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G29gat), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n437_), .A2(new_n439_), .A3(new_n431_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n435_), .A2(new_n440_), .A3(new_n428_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n427_), .B1(new_n434_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n432_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n428_), .B1(new_n435_), .B2(new_n440_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(KEYINPUT15), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT66), .ZN(new_n447_));
  OAI22_X1  g246(.A1(new_n447_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(KEYINPUT66), .B2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n447_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT65), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT65), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT6), .ZN(new_n455_));
  AND2_X1   g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n450_), .B(new_n451_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT8), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT67), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n465_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n459_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n460_), .A2(KEYINPUT9), .A3(new_n461_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT10), .B(G99gat), .ZN(new_n472_));
  OAI221_X1 g271(.A(new_n471_), .B1(KEYINPUT9), .B2(new_n461_), .C1(new_n472_), .C2(G106gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n457_), .A2(new_n458_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n469_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n426_), .B1(new_n446_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n424_), .A2(new_n425_), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n478_), .B(KEYINPUT72), .Z(new_n479_));
  INV_X1    g278(.A(KEYINPUT74), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n459_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n467_), .B1(new_n459_), .B2(new_n463_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n473_), .A2(new_n474_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n443_), .A2(new_n444_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n477_), .A2(new_n481_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n479_), .A2(new_n480_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n490_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G190gat), .B(G218gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(G134gat), .ZN(new_n495_));
  INV_X1    g294(.A(G162gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n497_), .B(new_n498_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n491_), .A2(new_n501_), .A3(new_n492_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT68), .B(G71gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(G78gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(G57gat), .B(G64gat), .Z(new_n506_));
  INV_X1    g305(.A(KEYINPUT11), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n507_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n505_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G78gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n504_), .B(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n508_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G231gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518_));
  INV_X1    g317(.A(G8gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G1gat), .B(G8gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n517_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT16), .B(G183gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G211gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G127gat), .B(G155gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  NOR3_X1   g328(.A1(new_n524_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(KEYINPUT17), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n524_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n422_), .A2(new_n503_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT12), .ZN(new_n535_));
  INV_X1    g334(.A(new_n515_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n476_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n537_), .B2(KEYINPUT69), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT69), .ZN(new_n539_));
  AOI211_X1 g338(.A(new_n539_), .B(KEYINPUT12), .C1(new_n476_), .C2(new_n536_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT70), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G230gat), .A2(G233gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT64), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n485_), .A2(new_n515_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n541_), .A2(new_n542_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT69), .B1(new_n485_), .B2(new_n515_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT12), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n537_), .A2(KEYINPUT69), .A3(new_n535_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n549_), .A2(new_n545_), .A3(new_n546_), .A4(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT70), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n545_), .B1(new_n546_), .B2(new_n537_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G120gat), .B(G148gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(new_n234_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT5), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n298_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n553_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT13), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n562_), .A2(new_n566_), .A3(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(new_n237_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT75), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n569_), .B(G197gat), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT75), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n571_), .A2(new_n574_), .A3(G169gat), .ZN(new_n575_));
  AOI21_X1  g374(.A(G169gat), .B1(new_n571_), .B2(new_n574_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n442_), .A2(new_n445_), .A3(new_n523_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n523_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n486_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n579_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n580_), .A2(new_n486_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n523_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n583_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n577_), .B1(new_n582_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n582_), .A2(new_n586_), .A3(new_n577_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT77), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n589_), .A2(KEYINPUT76), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n589_), .B2(KEYINPUT76), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n588_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(KEYINPUT76), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT77), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(KEYINPUT76), .A3(new_n590_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n587_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n568_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT102), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n534_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n202_), .B1(new_n601_), .B2(new_n384_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT103), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n593_), .A2(new_n597_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT78), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n422_), .A2(new_n605_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n503_), .A2(KEYINPUT37), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n503_), .A2(KEYINPUT37), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n533_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(new_n568_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n612_), .A2(G1gat), .A3(new_n383_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(KEYINPUT104), .B2(KEYINPUT38), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n615_));
  OAI211_X1 g414(.A(new_n603_), .B(new_n614_), .C1(new_n613_), .C2(new_n615_), .ZN(G1324gat));
  INV_X1    g415(.A(KEYINPUT105), .ZN(new_n617_));
  INV_X1    g416(.A(new_n354_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n534_), .A2(new_n617_), .A3(new_n618_), .A4(new_n600_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n396_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n284_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n278_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n384_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n623_), .A2(new_n354_), .B1(new_n418_), .B2(new_n285_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n394_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n620_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n533_), .A2(new_n503_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n600_), .A2(new_n626_), .A3(new_n618_), .A4(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT105), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n619_), .A2(new_n629_), .A3(G8gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT39), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n619_), .A2(new_n629_), .A3(new_n632_), .A4(G8gat), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n612_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n519_), .A3(new_n618_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(KEYINPUT40), .A3(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1325gat));
  INV_X1    g440(.A(G15gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n601_), .B2(new_n625_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT41), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n635_), .A2(new_n642_), .A3(new_n625_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1326gat));
  INV_X1    g445(.A(G22gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n621_), .A2(new_n622_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n635_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n601_), .A2(new_n648_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(G22gat), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT42), .B(new_n647_), .C1(new_n601_), .C2(new_n648_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT106), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(new_n649_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1327gat));
  INV_X1    g457(.A(new_n503_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n532_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n606_), .A2(new_n568_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G29gat), .B1(new_n662_), .B2(new_n384_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n600_), .A2(new_n533_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n609_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n666_), .B2(KEYINPUT107), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n626_), .B2(new_n609_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n625_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n609_), .B(new_n667_), .C1(new_n669_), .C2(new_n396_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n665_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(KEYINPUT108), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675_));
  INV_X1    g474(.A(new_n667_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n422_), .B2(new_n666_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n664_), .B1(new_n677_), .B2(new_n670_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n675_), .B1(new_n678_), .B2(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(new_n383_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n436_), .B1(new_n678_), .B2(KEYINPUT44), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n663_), .B1(new_n682_), .B2(new_n683_), .ZN(G1328gat));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n354_), .B1(new_n678_), .B2(KEYINPUT44), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n431_), .B1(new_n680_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n618_), .A2(new_n431_), .ZN(new_n689_));
  OR3_X1    g488(.A1(new_n661_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n661_), .B2(new_n689_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n685_), .B1(new_n687_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n692_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n678_), .A2(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n618_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n679_), .B2(new_n674_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT46), .B(new_n694_), .C1(new_n697_), .C2(new_n431_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n693_), .A2(new_n698_), .ZN(G1329gat));
  INV_X1    g498(.A(G43gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n678_), .B2(KEYINPUT44), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT108), .B1(new_n672_), .B2(new_n673_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n678_), .A2(new_n675_), .A3(KEYINPUT44), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n625_), .B(new_n701_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n700_), .B1(new_n661_), .B2(new_n394_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n704_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1330gat));
  AOI21_X1  g508(.A(G50gat), .B1(new_n662_), .B2(new_n648_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n681_), .A2(new_n285_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n695_), .A2(G50gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(G1331gat));
  INV_X1    g512(.A(new_n568_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n610_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n422_), .B1(KEYINPUT110), .B2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n716_), .B(new_n604_), .C1(KEYINPUT110), .C2(new_n715_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n384_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  OAI21_X1  g519(.A(G57gat), .B1(new_n383_), .B2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n534_), .A2(new_n714_), .A3(new_n605_), .ZN(new_n722_));
  INV_X1    g521(.A(G57gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(KEYINPUT111), .B2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n719_), .B1(new_n721_), .B2(new_n724_), .ZN(G1332gat));
  OAI21_X1  g524(.A(G64gat), .B1(new_n722_), .B2(new_n354_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT48), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n354_), .A2(G64gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n717_), .B2(new_n728_), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n722_), .B2(new_n394_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT49), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT49), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n732_), .B(G71gat), .C1(new_n722_), .C2(new_n394_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  OR3_X1    g533(.A1(new_n717_), .A2(G71gat), .A3(new_n394_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT112), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n734_), .A2(new_n738_), .A3(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n722_), .B2(new_n285_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n718_), .A2(new_n512_), .A3(new_n648_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1335gat));
  NOR2_X1   g543(.A1(new_n568_), .A2(new_n598_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n626_), .A2(new_n660_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n384_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n677_), .A2(new_n670_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n749_), .A2(new_n533_), .A3(new_n745_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n384_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n751_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g551(.A(G92gat), .B1(new_n747_), .B2(new_n618_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n750_), .A2(new_n618_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(G92gat), .ZN(G1337gat));
  OR2_X1    g554(.A1(new_n394_), .A2(new_n472_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT113), .B1(new_n746_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n750_), .A2(new_n625_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(G99gat), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(G1338gat));
  OR3_X1    g560(.A1(new_n746_), .A2(G106gat), .A3(new_n285_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n749_), .A2(new_n533_), .A3(new_n648_), .A4(new_n745_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G106gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G106gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT53), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n769_), .B(new_n762_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1339gat));
  AOI211_X1 g570(.A(new_n554_), .B(new_n561_), .C1(new_n547_), .C2(new_n552_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT116), .B1(new_n772_), .B2(new_n604_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n563_), .A2(new_n774_), .A3(new_n598_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n541_), .A2(new_n546_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n544_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n551_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n547_), .B2(new_n552_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n561_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(KEYINPUT56), .B(new_n561_), .C1(new_n780_), .C2(new_n782_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n776_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n578_), .A2(new_n583_), .A3(new_n581_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n579_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n789_), .B(new_n790_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n589_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n564_), .A2(new_n788_), .A3(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n560_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n795_), .B2(new_n772_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT118), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n659_), .B1(new_n787_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n785_), .A2(new_n786_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n792_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(new_n563_), .A3(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n803_), .A2(new_n804_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n802_), .A2(new_n563_), .A3(new_n807_), .A4(new_n805_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n609_), .A3(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT57), .B(new_n659_), .C1(new_n787_), .C2(new_n798_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n801_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n533_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n610_), .A2(new_n568_), .A3(new_n605_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(KEYINPUT115), .Z(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n815_), .B(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n814_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n285_), .A2(new_n384_), .A3(new_n354_), .A4(new_n625_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT120), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT59), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n827_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n358_), .B(new_n605_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n358_), .B1(new_n824_), .B2(new_n604_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT121), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1340gat));
  OAI21_X1  g631(.A(new_n366_), .B1(new_n568_), .B2(KEYINPUT60), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n825_), .B(new_n833_), .C1(KEYINPUT60), .C2(new_n366_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n568_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n366_), .ZN(G1341gat));
  AOI21_X1  g635(.A(G127gat), .B1(new_n825_), .B2(new_n532_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n533_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g638(.A(G134gat), .B1(new_n825_), .B2(new_n503_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n666_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g641(.A1(new_n285_), .A2(new_n383_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n821_), .A2(new_n354_), .A3(new_n394_), .A4(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n604_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n204_), .ZN(G1344gat));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n568_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(new_n205_), .ZN(G1345gat));
  NOR2_X1   g647(.A1(new_n844_), .A2(new_n533_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT61), .B(G155gat), .Z(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1346gat));
  NOR3_X1   g650(.A1(new_n844_), .A2(new_n496_), .A3(new_n666_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n496_), .B1(new_n844_), .B2(new_n659_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n853_), .A2(KEYINPUT122), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(KEYINPUT122), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n852_), .B1(new_n854_), .B2(new_n855_), .ZN(G1347gat));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n354_), .A2(new_n384_), .A3(new_n394_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n821_), .A2(new_n285_), .A3(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n604_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n857_), .B1(new_n860_), .B2(new_n297_), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT123), .B(G169gat), .C1(new_n859_), .C2(new_n604_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(KEYINPUT62), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n309_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n857_), .B(new_n865_), .C1(new_n860_), .C2(new_n297_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n864_), .A3(new_n866_), .ZN(G1348gat));
  NOR2_X1   g666(.A1(new_n859_), .A2(new_n568_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n298_), .ZN(G1349gat));
  NOR2_X1   g668(.A1(new_n859_), .A2(new_n533_), .ZN(new_n870_));
  MUX2_X1   g669(.A(G183gat), .B(new_n303_), .S(new_n870_), .Z(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n859_), .B2(new_n666_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n503_), .A2(new_n324_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n859_), .B2(new_n873_), .ZN(G1351gat));
  AOI21_X1  g673(.A(new_n819_), .B1(new_n813_), .B2(new_n533_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n623_), .A2(new_n394_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT124), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n875_), .A2(new_n354_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n598_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n714_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT125), .B(G204gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1353gat));
  AOI21_X1  g682(.A(new_n354_), .B1(new_n814_), .B2(new_n820_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n877_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT63), .B(G211gat), .Z(new_n886_));
  NAND4_X1  g685(.A1(new_n884_), .A2(new_n532_), .A3(new_n885_), .A4(new_n886_), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n875_), .A2(new_n533_), .A3(new_n354_), .A4(new_n877_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT126), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT127), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n887_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(new_n893_), .A3(new_n895_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n821_), .A2(new_n532_), .A3(new_n618_), .A4(new_n885_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n889_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n894_), .B1(new_n898_), .B2(new_n887_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n895_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT127), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n896_), .A2(new_n901_), .ZN(G1354gat));
  AOI21_X1  g701(.A(G218gat), .B1(new_n878_), .B2(new_n503_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n878_), .A2(new_n609_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(G218gat), .B2(new_n904_), .ZN(G1355gat));
endmodule


