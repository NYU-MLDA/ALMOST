//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT25), .B(G183gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n215_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n205_), .A2(new_n210_), .A3(new_n214_), .A4(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n208_), .B(new_n209_), .C1(G183gat), .C2(G190gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G227gat), .A2(G233gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(G15gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n223_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G71gat), .B(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G43gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT77), .B(KEYINPUT30), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n226_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n226_), .A2(new_n231_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT78), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G127gat), .B(G134gat), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(KEYINPUT79), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(KEYINPUT79), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G113gat), .B(G120gat), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT31), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n242_), .A2(KEYINPUT31), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n235_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n245_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(KEYINPUT80), .A3(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n234_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT78), .B1(new_n232_), .B2(new_n233_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n202_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n253_), .A2(KEYINPUT81), .A3(new_n234_), .A4(new_n249_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n232_), .A2(new_n233_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT84), .ZN(new_n261_));
  NOR3_X1   g060(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n269_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT1), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT82), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n277_), .A3(KEYINPUT1), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n273_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n280_));
  XOR2_X1   g079(.A(G141gat), .B(G148gat), .Z(new_n281_));
  AND3_X1   g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n280_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n259_), .B(new_n271_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT28), .B(G22gat), .ZN(new_n285_));
  INV_X1    g084(.A(G50gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n279_), .A2(new_n281_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT83), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n287_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n292_), .A2(new_n259_), .A3(new_n293_), .A4(new_n271_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n288_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n295_), .B1(new_n288_), .B2(new_n294_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT90), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n295_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n270_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n293_), .B1(new_n302_), .B2(new_n259_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n284_), .A2(new_n287_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n299_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT90), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n288_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G211gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(G218gat), .ZN(new_n310_));
  INV_X1    g109(.A(G218gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(G211gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT89), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT88), .ZN(new_n314_));
  INV_X1    g113(.A(G197gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(G204gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(G204gat), .ZN(new_n317_));
  INV_X1    g116(.A(G204gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n311_), .A2(G211gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n309_), .A2(G218gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n313_), .A2(new_n320_), .A3(KEYINPUT21), .A4(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n315_), .B2(G204gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n318_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n317_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n329_), .A2(KEYINPUT21), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT21), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n316_), .A2(new_n319_), .A3(new_n331_), .A4(new_n317_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n310_), .A2(new_n312_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n325_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n302_), .B2(new_n259_), .ZN(new_n336_));
  INV_X1    g135(.A(G228gat), .ZN(new_n337_));
  INV_X1    g136(.A(G233gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  OAI221_X1 g139(.A(new_n335_), .B1(new_n337_), .B2(new_n338_), .C1(new_n302_), .C2(new_n259_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n298_), .A2(new_n308_), .A3(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G78gat), .B(G106gat), .Z(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n341_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n345_), .B(KEYINPUT90), .C1(new_n296_), .C2(new_n297_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n343_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n344_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G1gat), .B(G29gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G57gat), .B(G85gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT94), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n271_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n302_), .A2(new_n242_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n357_), .A2(KEYINPUT4), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n357_), .B2(KEYINPUT4), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n355_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT4), .ZN(new_n365_));
  OR3_X1    g164(.A1(new_n302_), .A2(new_n242_), .A3(KEYINPUT4), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(KEYINPUT94), .A4(new_n361_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n354_), .B1(new_n364_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n354_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n363_), .A2(new_n368_), .A3(new_n371_), .A4(new_n367_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n349_), .A2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n220_), .A2(G169gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n211_), .A2(KEYINPUT22), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT91), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n211_), .A2(KEYINPUT22), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n220_), .A2(G169gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT91), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(G176gat), .B1(new_n377_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n218_), .A2(new_n215_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n217_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n335_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n329_), .A2(KEYINPUT21), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n387_), .A2(new_n222_), .A3(new_n217_), .A4(new_n325_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(KEYINPUT20), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n218_), .A2(new_n215_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n377_), .A2(new_n381_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(G176gat), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n395_), .A2(new_n217_), .A3(new_n387_), .A4(new_n325_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n391_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n335_), .A2(new_n223_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n396_), .A2(KEYINPUT20), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n392_), .A2(KEYINPUT92), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT92), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n389_), .A2(new_n401_), .A3(new_n391_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT18), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT27), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n398_), .B(KEYINPUT20), .C1(new_n335_), .C2(new_n384_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n391_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n391_), .B2(new_n389_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n410_), .B1(new_n413_), .B2(new_n407_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n384_), .B2(new_n335_), .ZN(new_n417_));
  AOI211_X1 g216(.A(KEYINPUT92), .B(new_n397_), .C1(new_n417_), .C2(new_n388_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n401_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n399_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT93), .B1(new_n420_), .B2(new_n407_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT93), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n403_), .A2(new_n422_), .A3(new_n408_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n400_), .A2(new_n407_), .A3(new_n402_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n415_), .B1(new_n425_), .B2(new_n410_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n374_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n407_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n428_), .B2(new_n422_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n420_), .A2(KEYINPUT93), .A3(new_n407_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n357_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n354_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n366_), .A2(new_n360_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n365_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n372_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n369_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n438_), .A2(KEYINPUT33), .A3(new_n371_), .A4(new_n363_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n431_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n408_), .A2(KEYINPUT32), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n420_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n441_), .B2(new_n413_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n373_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n349_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n258_), .B1(new_n427_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n373_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n258_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT96), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n349_), .A2(new_n451_), .A3(new_n426_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n349_), .B2(new_n426_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n450_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT97), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n410_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n343_), .A2(new_n346_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n344_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n343_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n409_), .A2(new_n414_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n457_), .A2(new_n460_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT96), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n349_), .A2(new_n426_), .A3(new_n451_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(KEYINPUT97), .A3(new_n450_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n447_), .B1(new_n456_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G113gat), .B(G141gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G169gat), .B(G197gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n469_), .B(new_n470_), .Z(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT76), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT74), .B(G1gat), .ZN(new_n474_));
  INV_X1    g273(.A(G8gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT75), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G1gat), .B(G8gat), .Z(new_n480_));
  AND2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n479_), .A2(new_n480_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G29gat), .B(G36gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G43gat), .B(G50gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n473_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(KEYINPUT76), .B(new_n486_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n488_), .A2(new_n489_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G229gat), .A2(G233gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n489_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n486_), .B(KEYINPUT15), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n483_), .A2(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n493_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n472_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n488_), .A2(new_n489_), .B1(new_n483_), .B2(new_n494_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n491_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n499_), .B(new_n471_), .C1(new_n491_), .C2(new_n490_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n468_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT66), .ZN(new_n505_));
  XOR2_X1   g304(.A(G85gat), .B(G92gat), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT9), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT64), .B(G92gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT9), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(G85gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT65), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT6), .Z(new_n514_));
  INV_X1    g313(.A(G106gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT7), .Z(new_n520_));
  OAI21_X1  g319(.A(new_n506_), .B1(new_n520_), .B2(new_n514_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT8), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n526_));
  XOR2_X1   g325(.A(G71gat), .B(G78gat), .Z(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n526_), .A2(new_n527_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n505_), .B1(new_n523_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n504_), .A2(KEYINPUT66), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n523_), .A2(new_n531_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n523_), .B2(new_n531_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n533_), .B(new_n534_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n534_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n518_), .A2(new_n522_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(new_n530_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n523_), .A2(new_n531_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n541_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G120gat), .B(G148gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT5), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G176gat), .B(G204gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(KEYINPUT67), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT68), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n546_), .B(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT13), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(KEYINPUT13), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n523_), .A2(new_n494_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT34), .ZN(new_n560_));
  OAI221_X1 g359(.A(new_n558_), .B1(KEYINPUT35), .B2(new_n560_), .C1(new_n487_), .C2(new_n523_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n560_), .A2(KEYINPUT35), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n562_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT69), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT36), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT70), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(KEYINPUT71), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n565_), .A2(new_n572_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT71), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n569_), .B(KEYINPUT36), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n565_), .A2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(KEYINPUT37), .B(new_n573_), .C1(new_n576_), .C2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n563_), .A2(new_n564_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT72), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n578_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n582_), .B2(new_n581_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n574_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n580_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n530_), .B(new_n589_), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n483_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593_));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT16), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  OR3_X1    g396(.A1(new_n592_), .A2(new_n593_), .A3(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(KEYINPUT17), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n592_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n588_), .A2(new_n601_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n503_), .A2(new_n557_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n373_), .A3(new_n474_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT38), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n584_), .A2(new_n574_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n468_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n557_), .A2(new_n501_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n601_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n448_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n604_), .A2(new_n605_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n606_), .A2(new_n614_), .A3(new_n615_), .ZN(G1324gat));
  INV_X1    g415(.A(new_n426_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n612_), .A2(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n618_), .A2(KEYINPUT98), .A3(G8gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT98), .B1(new_n618_), .B2(G8gat), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n621_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n603_), .A2(new_n475_), .A3(new_n617_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT40), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT40), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(G1325gat));
  INV_X1    g429(.A(G15gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n612_), .B2(new_n258_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT41), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n603_), .A2(new_n631_), .A3(new_n258_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(G1326gat));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n349_), .B(KEYINPUT99), .Z(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n612_), .B2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n603_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1327gat));
  INV_X1    g441(.A(new_n601_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n607_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(new_n557_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n503_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G29gat), .B1(new_n647_), .B2(new_n373_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n610_), .A2(new_n643_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n468_), .A2(KEYINPUT43), .A3(new_n587_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n427_), .A2(new_n446_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n258_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT97), .B1(new_n466_), .B2(new_n450_), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n455_), .B(new_n449_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n654_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n651_), .B1(new_n657_), .B2(new_n588_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n649_), .B1(new_n650_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT44), .B(new_n649_), .C1(new_n650_), .C2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n373_), .A2(G29gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n648_), .B1(new_n664_), .B2(new_n665_), .ZN(G1328gat));
  OR2_X1    g465(.A1(new_n426_), .A2(KEYINPUT102), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n426_), .A2(KEYINPUT102), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n646_), .A2(G36gat), .A3(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT45), .Z(new_n672_));
  NAND3_X1  g471(.A1(new_n661_), .A2(new_n617_), .A3(new_n662_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n673_), .A2(new_n674_), .A3(G36gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n673_), .B2(G36gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT46), .B(new_n672_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  OAI21_X1  g480(.A(new_n228_), .B1(new_n646_), .B2(new_n653_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n258_), .A2(G43gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n663_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686_));
  INV_X1    g485(.A(new_n349_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n664_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G50gat), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n647_), .A2(new_n286_), .A3(new_n637_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n686_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT103), .B(new_n690_), .C1(new_n688_), .C2(G50gat), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1331gat));
  NOR3_X1   g493(.A1(new_n557_), .A2(new_n501_), .A3(new_n601_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n609_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G57gat), .B1(new_n697_), .B2(new_n448_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n557_), .A2(new_n501_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n657_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(new_n602_), .ZN(new_n701_));
  INV_X1    g500(.A(G57gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n373_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n698_), .A2(new_n703_), .ZN(G1332gat));
  INV_X1    g503(.A(G64gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n696_), .B2(new_n669_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT48), .Z(new_n707_));
  NAND3_X1  g506(.A1(new_n701_), .A2(new_n705_), .A3(new_n669_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n707_), .A2(KEYINPUT104), .A3(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1333gat));
  INV_X1    g512(.A(G71gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n696_), .B2(new_n258_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT49), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n701_), .A2(new_n714_), .A3(new_n258_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1334gat));
  INV_X1    g517(.A(G78gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n696_), .B2(new_n637_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT50), .Z(new_n721_));
  NAND3_X1  g520(.A1(new_n701_), .A2(new_n719_), .A3(new_n637_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1335gat));
  NAND2_X1  g522(.A1(new_n699_), .A2(new_n601_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT43), .B1(new_n468_), .B2(new_n587_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n657_), .A2(new_n651_), .A3(new_n588_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G85gat), .B1(new_n728_), .B2(new_n448_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n700_), .A2(new_n644_), .ZN(new_n730_));
  INV_X1    g529(.A(G85gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n373_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n729_), .A2(new_n732_), .ZN(G1336gat));
  AOI21_X1  g532(.A(G92gat), .B1(new_n730_), .B2(new_n617_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT105), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n669_), .A2(new_n508_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n727_), .B2(new_n736_), .ZN(G1337gat));
  OAI21_X1  g536(.A(G99gat), .B1(new_n728_), .B2(new_n653_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n730_), .A2(new_n258_), .A3(new_n516_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g541(.A1(new_n730_), .A2(new_n515_), .A3(new_n687_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744_));
  INV_X1    g543(.A(new_n724_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n687_), .B(new_n745_), .C1(new_n650_), .C2(new_n658_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G106gat), .B1(new_n746_), .B2(KEYINPUT107), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n727_), .B2(new_n687_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n744_), .B1(new_n748_), .B2(new_n751_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n747_), .A2(new_n750_), .A3(KEYINPUT52), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n743_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n743_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1339gat));
  INV_X1    g557(.A(KEYINPUT118), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n587_), .A2(new_n502_), .A3(new_n557_), .A4(new_n643_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n761_), .A2(KEYINPUT54), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(KEYINPUT54), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT109), .Z(new_n764_));
  AND3_X1   g563(.A1(new_n760_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n760_), .B2(new_n762_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n535_), .B1(new_n542_), .B2(new_n530_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n532_), .B1(new_n769_), .B2(new_n537_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n770_), .A2(new_n534_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n770_), .B2(new_n534_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n540_), .A2(KEYINPUT110), .A3(new_n774_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT56), .B(new_n550_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT114), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n774_), .B1(new_n540_), .B2(KEYINPUT110), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n773_), .A2(new_n774_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n771_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(KEYINPUT56), .A4(new_n550_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n770_), .A2(new_n534_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n776_), .A2(new_n779_), .A3(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n787_), .B2(new_n551_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n778_), .A2(new_n784_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(KEYINPUT58), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n540_), .A2(new_n545_), .A3(new_n551_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n491_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n472_), .B1(new_n490_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n493_), .A2(new_n495_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n491_), .B1(new_n797_), .B2(KEYINPUT111), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n498_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n796_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n492_), .A2(new_n496_), .A3(new_n472_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT112), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n804_));
  INV_X1    g603(.A(new_n800_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n795_), .B1(new_n498_), .B2(new_n799_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n804_), .B(new_n500_), .C1(new_n807_), .C2(new_n796_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n794_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n789_), .A2(new_n792_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n792_), .B1(new_n789_), .B2(new_n809_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n810_), .A2(new_n811_), .A3(new_n587_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n501_), .A2(new_n793_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n788_), .B2(new_n777_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n554_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n607_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n768_), .B1(new_n812_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n789_), .A2(new_n809_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n791_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n789_), .A2(new_n809_), .A3(new_n792_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n588_), .A3(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT117), .A3(new_n819_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n817_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT57), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n821_), .A2(new_n826_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n767_), .B1(new_n829_), .B2(new_n601_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n466_), .A2(new_n258_), .A3(new_n373_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n831_), .A2(KEYINPUT116), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(KEYINPUT116), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n759_), .B1(new_n830_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n835_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n825_), .A2(new_n819_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n838_), .A2(new_n768_), .B1(KEYINPUT57), .B2(new_n827_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n643_), .B1(new_n839_), .B2(new_n826_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT118), .B(new_n837_), .C1(new_n840_), .C2(new_n767_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n819_), .A2(KEYINPUT113), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n817_), .A2(new_n843_), .A3(new_n818_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n842_), .A2(new_n825_), .A3(new_n828_), .A4(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n767_), .B1(new_n601_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT59), .B1(new_n846_), .B2(new_n831_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n836_), .A2(new_n841_), .A3(new_n501_), .A4(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G113gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n846_), .A2(new_n831_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  OR3_X1    g650(.A1(new_n851_), .A2(G113gat), .A3(new_n502_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n852_), .ZN(G1340gat));
  INV_X1    g652(.A(new_n557_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n836_), .A2(new_n841_), .A3(new_n854_), .A4(new_n847_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G120gat), .ZN(new_n856_));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n557_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT119), .B1(new_n857_), .B2(KEYINPUT60), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n850_), .B(new_n860_), .C1(new_n861_), .C2(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n856_), .A2(new_n862_), .ZN(G1341gat));
  NAND4_X1  g662(.A1(new_n836_), .A2(new_n841_), .A3(new_n643_), .A4(new_n847_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G127gat), .ZN(new_n865_));
  OR3_X1    g664(.A1(new_n851_), .A2(G127gat), .A3(new_n601_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1342gat));
  NAND4_X1  g666(.A1(new_n836_), .A2(new_n841_), .A3(new_n588_), .A4(new_n847_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G134gat), .ZN(new_n869_));
  OR3_X1    g668(.A1(new_n851_), .A2(G134gat), .A3(new_n607_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1343gat));
  NOR3_X1   g670(.A1(new_n669_), .A2(new_n349_), .A3(new_n448_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n846_), .A2(new_n258_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n501_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n854_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n643_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1346gat));
  NAND2_X1  g680(.A1(new_n874_), .A2(new_n608_), .ZN(new_n882_));
  INV_X1    g681(.A(G162gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(KEYINPUT120), .A3(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885_));
  NOR4_X1   g684(.A1(new_n846_), .A2(new_n258_), .A3(new_n607_), .A4(new_n873_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(G162gat), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n587_), .A2(new_n883_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n884_), .A2(new_n887_), .B1(new_n874_), .B2(new_n888_), .ZN(G1347gat));
  NAND2_X1  g688(.A1(new_n669_), .A2(new_n450_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n637_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n501_), .B(new_n891_), .C1(new_n840_), .C2(new_n767_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G169gat), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n894_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n892_), .A2(G169gat), .A3(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n895_), .B(new_n897_), .C1(new_n394_), .C2(new_n892_), .ZN(G1348gat));
  INV_X1    g697(.A(new_n891_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n830_), .A2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G176gat), .B1(new_n900_), .B2(new_n854_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n846_), .A2(new_n687_), .A3(new_n890_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n557_), .A2(new_n212_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(KEYINPUT122), .A3(new_n903_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n901_), .B1(new_n906_), .B2(new_n907_), .ZN(G1349gat));
  AOI21_X1  g707(.A(G183gat), .B1(new_n902_), .B2(new_n643_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n601_), .A2(new_n203_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n900_), .B2(new_n910_), .ZN(G1350gat));
  NAND3_X1  g710(.A1(new_n900_), .A2(new_n204_), .A3(new_n608_), .ZN(new_n912_));
  INV_X1    g711(.A(G190gat), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n830_), .A2(new_n587_), .A3(new_n899_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1351gat));
  NOR2_X1   g714(.A1(new_n846_), .A2(new_n258_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n669_), .A2(new_n374_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(new_n501_), .A3(new_n918_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n315_), .A2(KEYINPUT123), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT123), .B(G197gat), .Z(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n919_), .B2(new_n922_), .ZN(G1352gat));
  NAND3_X1  g722(.A1(new_n916_), .A2(new_n854_), .A3(new_n918_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g724(.A(new_n601_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT124), .Z(new_n927_));
  NAND3_X1  g726(.A1(new_n916_), .A2(new_n918_), .A3(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n929_));
  NOR3_X1   g728(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT126), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n928_), .A2(new_n929_), .A3(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1354gat));
  NOR2_X1   g733(.A1(new_n607_), .A2(G218gat), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n916_), .A2(new_n918_), .A3(new_n935_), .ZN(new_n936_));
  NOR4_X1   g735(.A1(new_n846_), .A2(new_n258_), .A3(new_n587_), .A4(new_n917_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(new_n311_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(KEYINPUT127), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n936_), .B(new_n940_), .C1(new_n937_), .C2(new_n311_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1355gat));
endmodule


