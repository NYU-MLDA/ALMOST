//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G155gat), .B(G162gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n208_), .B(KEYINPUT87), .C1(KEYINPUT1), .C2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT87), .ZN(new_n211_));
  AND2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NOR3_X1   g012(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT1), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n211_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n209_), .A2(KEYINPUT88), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n205_), .A2(KEYINPUT3), .ZN(new_n219_));
  OR3_X1    g018(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n207_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n219_), .A2(new_n220_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n209_), .A2(KEYINPUT88), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n218_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G127gat), .B(G134gat), .Z(new_n227_));
  XOR2_X1   g026(.A(G113gat), .B(G120gat), .Z(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n217_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n217_), .B2(new_n226_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT93), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n217_), .A2(new_n226_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n229_), .ZN(new_n235_));
  NOR3_X1   g034(.A1(new_n234_), .A2(KEYINPUT93), .A3(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n202_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n235_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n217_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT93), .A3(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n217_), .A2(new_n226_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(new_n232_), .A3(new_n229_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n238_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n231_), .A2(new_n238_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n202_), .B(KEYINPUT94), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n237_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G1gat), .B(G29gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G85gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT0), .B(G57gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n250_), .B(new_n251_), .Z(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n237_), .B(new_n252_), .C1(new_n244_), .C2(new_n247_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT29), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n242_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n234_), .B2(KEYINPUT29), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(G228gat), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G78gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G106gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n263_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G197gat), .A2(G204gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT91), .B(G204gat), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(G197gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G211gat), .B(G218gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT21), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n274_), .A2(KEYINPUT21), .ZN(new_n279_));
  OR2_X1    g078(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n280_));
  INV_X1    g079(.A(G197gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n276_), .B1(G197gat), .B2(G204gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n275_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n278_), .B1(new_n279_), .B2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G22gat), .B(G50gat), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n287_), .B(new_n289_), .C1(new_n242_), .C2(new_n258_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n258_), .B1(new_n217_), .B2(new_n226_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n287_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n288_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n270_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n261_), .A2(new_n294_), .A3(new_n262_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n271_), .A2(new_n290_), .A3(new_n293_), .A4(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n293_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n261_), .A2(new_n294_), .A3(new_n262_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n294_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT20), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT23), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(G183gat), .B2(G190gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(G169gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT25), .B(G183gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT26), .B(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT24), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(G169gat), .B2(G176gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(G169gat), .B2(G176gat), .ZN(new_n314_));
  OR3_X1    g113(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n311_), .A2(new_n314_), .A3(new_n304_), .A4(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n308_), .A2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n302_), .B1(new_n317_), .B2(new_n287_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n304_), .A2(new_n315_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT83), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n321_));
  NAND2_X1  g120(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT26), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n325_));
  INV_X1    g124(.A(G183gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n323_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(G183gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(G183gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n330_), .B1(new_n331_), .B2(KEYINPUT80), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n314_), .B(new_n321_), .C1(new_n328_), .C2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT83), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n304_), .A2(new_n334_), .A3(new_n315_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n320_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n314_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n337_), .A2(KEYINPUT82), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n308_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n318_), .B1(new_n339_), .B2(new_n287_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G226gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT19), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G8gat), .B(G36gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n339_), .A2(new_n287_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n342_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n308_), .A2(new_n316_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n302_), .B1(new_n292_), .B2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n343_), .A2(new_n349_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n343_), .A2(new_n354_), .A3(KEYINPUT96), .A4(new_n349_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n318_), .B(new_n351_), .C1(new_n339_), .C2(new_n287_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT20), .B1(new_n317_), .B2(new_n287_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n339_), .B2(new_n287_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n359_), .B1(new_n361_), .B2(new_n351_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n348_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n357_), .A2(new_n358_), .A3(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n364_), .A2(KEYINPUT27), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n343_), .A2(new_n349_), .A3(new_n354_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n349_), .B1(new_n343_), .B2(new_n354_), .ZN(new_n367_));
  OR3_X1    g166(.A1(new_n366_), .A2(new_n367_), .A3(KEYINPUT27), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n257_), .B(new_n301_), .C1(new_n365_), .C2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT33), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n255_), .A2(KEYINPUT95), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT95), .B1(new_n255_), .B2(new_n371_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n366_), .A2(new_n367_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n246_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n245_), .A2(new_n202_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n376_), .B(new_n253_), .C1(new_n244_), .C2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n255_), .B2(new_n371_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n362_), .A2(KEYINPUT32), .A3(new_n349_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n343_), .A2(new_n354_), .A3(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n374_), .A2(new_n380_), .B1(new_n256_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n370_), .B1(new_n385_), .B2(new_n301_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT84), .B(G43gat), .ZN(new_n388_));
  INV_X1    g187(.A(G99gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT30), .B(new_n308_), .C1(new_n336_), .C2(new_n338_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n337_), .A2(KEYINPUT82), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n394_), .A2(new_n333_), .A3(new_n320_), .A4(new_n335_), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT30), .B1(new_n395_), .B2(new_n308_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(G15gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(G71gat), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n393_), .A2(new_n396_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n339_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n404_), .B2(new_n392_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n391_), .B1(new_n401_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n400_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n392_), .A3(new_n402_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n390_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n387_), .B1(new_n410_), .B2(KEYINPUT85), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412_));
  AOI211_X1 g211(.A(new_n412_), .B(KEYINPUT86), .C1(new_n406_), .C2(new_n409_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n410_), .A2(KEYINPUT85), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n229_), .B(KEYINPUT31), .ZN(new_n415_));
  OAI22_X1  g214(.A1(new_n411_), .A2(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n407_), .A2(new_n390_), .A3(new_n408_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n390_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n419_), .B2(new_n412_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT85), .B1(new_n417_), .B2(new_n418_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT86), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n410_), .A2(KEYINPUT85), .A3(new_n387_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n416_), .A2(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n416_), .A2(new_n424_), .A3(new_n257_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n364_), .A2(KEYINPUT27), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n301_), .B1(new_n427_), .B2(new_n368_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n386_), .A2(new_n425_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G113gat), .B(G141gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G169gat), .B(G197gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n430_), .B(new_n431_), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G29gat), .B(G36gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT74), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G43gat), .B(G50gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT15), .ZN(new_n438_));
  INV_X1    g237(.A(new_n436_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n435_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT15), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT77), .B(G8gat), .ZN(new_n444_));
  INV_X1    g243(.A(G1gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT14), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G15gat), .B(G22gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT78), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G1gat), .B(G8gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n448_), .B(KEYINPUT78), .ZN(new_n453_));
  INV_X1    g252(.A(new_n451_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n443_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n455_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n437_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G229gat), .A2(G233gat), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n456_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n452_), .A2(new_n455_), .A3(new_n440_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n433_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n462_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n456_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n432_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n429_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT13), .ZN(new_n470_));
  XOR2_X1   g269(.A(KEYINPUT10), .B(G99gat), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n269_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G85gat), .B(G92gat), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT9), .ZN(new_n474_));
  INV_X1    g273(.A(G85gat), .ZN(new_n475_));
  INV_X1    g274(.A(G92gat), .ZN(new_n476_));
  OR3_X1    g275(.A1(new_n475_), .A2(new_n476_), .A3(KEYINPUT9), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT6), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n472_), .A2(new_n474_), .A3(new_n477_), .A4(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n389_), .A2(new_n269_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n479_), .A2(new_n481_), .B1(new_n484_), .B2(KEYINPUT7), .ZN(new_n485_));
  NAND2_X1  g284(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(new_n389_), .A3(new_n269_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT65), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n488_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT65), .ZN(new_n491_));
  NOR2_X1   g290(.A1(G99gat), .A2(G106gat), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .A4(new_n486_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n485_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n495_));
  NAND2_X1  g294(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n473_), .A2(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n483_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT69), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT69), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(new_n483_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n505_));
  XOR2_X1   g304(.A(G71gat), .B(G78gat), .Z(new_n506_));
  OR2_X1    g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n506_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT12), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n501_), .A2(new_n503_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n500_), .A2(new_n511_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT12), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AND2_X1   g316(.A1(G230gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n483_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n494_), .A2(new_n497_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n495_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n519_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n518_), .B1(new_n524_), .B2(new_n510_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n514_), .A2(new_n517_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT70), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n514_), .A2(new_n517_), .A3(new_n528_), .A4(new_n525_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT68), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(KEYINPUT67), .A3(new_n510_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n483_), .B(new_n510_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n532_), .A2(new_n535_), .A3(new_n515_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n531_), .B1(new_n536_), .B2(new_n518_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n531_), .A3(new_n518_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G120gat), .B(G148gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT5), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G176gat), .B(G204gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n530_), .A2(new_n540_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n530_), .B2(new_n540_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n470_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n539_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n527_), .B(new_n529_), .C1(new_n550_), .C2(new_n537_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n544_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(new_n546_), .A3(KEYINPUT13), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT71), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(KEYINPUT73), .B(KEYINPUT35), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT75), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n565_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT75), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n443_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n563_), .A2(new_n564_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n524_), .B2(new_n437_), .ZN(new_n572_));
  AOI211_X1 g371(.A(new_n567_), .B(new_n569_), .C1(new_n570_), .C2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n570_), .A2(KEYINPUT75), .A3(new_n568_), .A4(new_n572_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n560_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n570_), .A2(new_n572_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n567_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n569_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n560_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n574_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n559_), .B1(new_n576_), .B2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n581_), .B1(new_n580_), .B2(new_n574_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT37), .B1(new_n584_), .B2(KEYINPUT76), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n583_), .B(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n510_), .B(new_n587_), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(new_n457_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G127gat), .B(G155gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT16), .ZN(new_n592_));
  XOR2_X1   g391(.A(G183gat), .B(G211gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n589_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n590_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OR3_X1    g396(.A1(new_n589_), .A2(KEYINPUT79), .A3(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n589_), .B2(KEYINPUT79), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n595_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n586_), .A2(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n469_), .A2(new_n555_), .A3(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n445_), .A3(new_n256_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT97), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT38), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n554_), .B2(new_n468_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n549_), .A2(KEYINPUT98), .A3(new_n467_), .A4(new_n553_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n611_), .B2(new_n600_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n583_), .B(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n429_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n600_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n609_), .A2(KEYINPUT99), .A3(new_n610_), .A4(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n615_), .A3(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n618_), .B2(new_n257_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n604_), .A2(new_n605_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n606_), .A2(new_n619_), .A3(new_n620_), .ZN(G1324gat));
  NOR2_X1   g420(.A1(new_n365_), .A2(new_n369_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n602_), .A2(new_n444_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n625_), .A2(new_n626_), .A3(G8gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n625_), .B2(G8gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n623_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g429(.A(new_n425_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n602_), .A2(new_n398_), .A3(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G15gat), .B1(new_n618_), .B2(new_n425_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(new_n634_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n635_), .B2(new_n636_), .ZN(G1326gat));
  INV_X1    g436(.A(G22gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n301_), .B(KEYINPUT101), .Z(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n602_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G22gat), .B1(new_n618_), .B2(new_n639_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n642_), .A2(KEYINPUT103), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(KEYINPUT103), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n641_), .B1(new_n646_), .B2(new_n647_), .ZN(G1327gat));
  NAND2_X1  g447(.A1(new_n614_), .A2(new_n600_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n554_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n469_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G29gat), .B1(new_n651_), .B2(new_n256_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n609_), .A2(new_n610_), .A3(new_n600_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n428_), .A2(new_n416_), .A3(new_n424_), .A4(new_n257_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n301_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n427_), .B2(new_n368_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n384_), .A2(new_n256_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n255_), .A2(new_n371_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n255_), .A2(KEYINPUT95), .A3(new_n371_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n366_), .A2(new_n367_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n663_), .B(new_n378_), .C1(new_n371_), .C2(new_n255_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n657_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n301_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n656_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n654_), .B1(new_n667_), .B2(new_n631_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n586_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n668_), .B2(new_n586_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n653_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n586_), .ZN(new_n675_));
  OAI21_X1  g474(.A(KEYINPUT43), .B1(new_n429_), .B2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n668_), .A2(new_n669_), .A3(new_n586_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n678_), .A2(KEYINPUT104), .A3(new_n653_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n674_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n653_), .B(KEYINPUT44), .C1(new_n670_), .C2(new_n671_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n256_), .A2(G29gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n652_), .B1(new_n683_), .B2(new_n684_), .ZN(G1328gat));
  INV_X1    g484(.A(new_n651_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n686_), .A2(G36gat), .A3(new_n624_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n683_), .A2(new_n622_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(G36gat), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT46), .ZN(G1329gat));
  NOR3_X1   g491(.A1(new_n686_), .A2(G43gat), .A3(new_n425_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n683_), .A2(new_n631_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G43gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g495(.A(G50gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n651_), .A2(new_n697_), .A3(new_n640_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n682_), .A2(new_n301_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT44), .B1(new_n672_), .B2(new_n673_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n679_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n701_), .B2(KEYINPUT106), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n609_), .A2(new_n610_), .A3(new_n600_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n666_), .B1(new_n704_), .B2(KEYINPUT44), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT106), .B1(new_n681_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT107), .B1(new_n702_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n680_), .B1(new_n704_), .B2(KEYINPUT104), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n672_), .A2(new_n673_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT106), .B(new_n705_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G50gat), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n712_), .A2(new_n713_), .A3(new_n706_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n698_), .B1(new_n708_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(KEYINPUT108), .B(new_n698_), .C1(new_n708_), .C2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1331gat));
  INV_X1    g518(.A(new_n555_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n600_), .A2(new_n467_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n615_), .A3(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT110), .ZN(new_n723_));
  OAI21_X1  g522(.A(G57gat), .B1(new_n257_), .B2(KEYINPUT111), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n723_), .B(new_n724_), .C1(KEYINPUT111), .C2(G57gat), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n429_), .A2(new_n467_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n554_), .A3(new_n601_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT109), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(new_n257_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(G57gat), .B2(new_n729_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT112), .Z(G1332gat));
  INV_X1    g530(.A(G64gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n723_), .B2(new_n622_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT48), .Z(new_n734_));
  INV_X1    g533(.A(new_n728_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n732_), .A3(new_n622_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n723_), .B2(new_n631_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT49), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n738_), .A3(new_n631_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1334gat));
  AOI21_X1  g541(.A(new_n267_), .B1(new_n723_), .B2(new_n640_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT50), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n735_), .A2(new_n267_), .A3(new_n640_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1335gat));
  NAND4_X1  g545(.A1(new_n678_), .A2(new_n468_), .A3(new_n554_), .A4(new_n600_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n257_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n720_), .A2(new_n726_), .A3(new_n600_), .A4(new_n614_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n475_), .A3(new_n256_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1336gat));
  OAI21_X1  g551(.A(G92gat), .B1(new_n747_), .B2(new_n624_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n476_), .A3(new_n622_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1337gat));
  OAI21_X1  g554(.A(G99gat), .B1(new_n747_), .B2(new_n425_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT113), .Z(new_n757_));
  NAND3_X1  g556(.A1(new_n750_), .A2(new_n471_), .A3(new_n631_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g559(.A(G106gat), .B1(new_n747_), .B2(new_n666_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT52), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n750_), .A2(new_n269_), .A3(new_n301_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g564(.A1(new_n631_), .A2(new_n256_), .A3(new_n428_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n458_), .A2(new_n461_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n459_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n456_), .A2(G229gat), .A3(new_n458_), .A4(G233gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n433_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n466_), .A2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n547_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n514_), .A2(new_n517_), .A3(new_n535_), .A4(new_n532_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n532_), .A2(new_n535_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n777_), .A2(KEYINPUT117), .A3(new_n514_), .A4(new_n517_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n518_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n527_), .A2(new_n781_), .A3(new_n529_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n526_), .A2(new_n781_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT56), .B1(new_n784_), .B2(new_n544_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(KEYINPUT56), .A3(new_n544_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(KEYINPUT118), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n784_), .A2(new_n788_), .A3(KEYINPUT56), .A4(new_n544_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n773_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n586_), .B1(new_n790_), .B2(KEYINPUT58), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n786_), .A2(KEYINPUT118), .ZN(new_n793_));
  INV_X1    g592(.A(new_n785_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n789_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n772_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n792_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n790_), .A2(KEYINPUT119), .A3(KEYINPUT58), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n791_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT116), .B1(new_n547_), .B2(new_n468_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n546_), .A2(new_n802_), .A3(new_n467_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n786_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n801_), .B(new_n803_), .C1(new_n804_), .C2(new_n785_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n771_), .B1(new_n552_), .B2(new_n546_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n614_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n809_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n614_), .B(new_n814_), .C1(new_n805_), .C2(new_n807_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n810_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n600_), .B1(new_n800_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n818_));
  OR2_X1    g617(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n549_), .A2(new_n553_), .A3(new_n721_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n586_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT115), .B(new_n819_), .C1(new_n820_), .C2(new_n586_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n823_), .A2(KEYINPUT114), .A3(KEYINPUT54), .A4(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n817_), .A2(new_n818_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n675_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT119), .B1(new_n790_), .B2(KEYINPUT58), .ZN(new_n833_));
  AND4_X1   g632(.A1(KEYINPUT119), .A2(new_n795_), .A3(KEYINPUT58), .A4(new_n772_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n805_), .A2(new_n807_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n614_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n813_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n616_), .B1(new_n835_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT121), .B1(new_n840_), .B2(new_n829_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n766_), .B1(new_n831_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n467_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n766_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n846_));
  OAI211_X1 g645(.A(new_n845_), .B(new_n846_), .C1(new_n840_), .C2(new_n829_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n467_), .B(new_n847_), .C1(new_n842_), .C2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n844_), .B1(new_n850_), .B2(new_n843_), .ZN(G1340gat));
  OAI21_X1  g650(.A(new_n847_), .B1(new_n842_), .B2(new_n848_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G120gat), .B1(new_n852_), .B2(new_n555_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n842_), .ZN(new_n854_));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  INV_X1    g654(.A(new_n554_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(KEYINPUT60), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(KEYINPUT60), .B2(new_n855_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n853_), .B1(new_n854_), .B2(new_n858_), .ZN(G1341gat));
  NAND2_X1  g658(.A1(new_n616_), .A2(G127gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT123), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n847_), .B(new_n861_), .C1(new_n842_), .C2(new_n848_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(G127gat), .B1(new_n842_), .B2(new_n616_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1342gat));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n842_), .A2(new_n866_), .A3(new_n614_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n586_), .B(new_n847_), .C1(new_n842_), .C2(new_n848_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n869_), .B2(new_n866_), .ZN(G1343gat));
  NAND2_X1  g669(.A1(new_n831_), .A2(new_n841_), .ZN(new_n871_));
  NOR4_X1   g670(.A1(new_n631_), .A2(new_n257_), .A3(new_n666_), .A4(new_n622_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n468_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n203_), .ZN(G1344gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n555_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n204_), .ZN(G1345gat));
  AOI21_X1  g676(.A(new_n818_), .B1(new_n817_), .B2(new_n830_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n840_), .A2(KEYINPUT121), .A3(new_n829_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n616_), .B(new_n872_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT124), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n871_), .A2(new_n882_), .A3(new_n616_), .A4(new_n872_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n881_), .A2(new_n883_), .A3(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n873_), .B2(new_n675_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n837_), .A2(G162gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n873_), .B2(new_n889_), .ZN(G1347gat));
  AOI21_X1  g689(.A(new_n640_), .B1(new_n817_), .B2(new_n830_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n624_), .A2(new_n425_), .A3(new_n256_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT22), .B(G169gat), .Z(new_n894_));
  NOR2_X1   g693(.A1(new_n468_), .A2(new_n894_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(KEYINPUT125), .Z(new_n896_));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n893_), .A2(new_n467_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(G169gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(G169gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n897_), .B1(new_n900_), .B2(new_n901_), .ZN(G1348gat));
  AOI21_X1  g701(.A(G176gat), .B1(new_n893_), .B2(new_n554_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n301_), .B1(new_n831_), .B2(new_n841_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n720_), .A2(G176gat), .A3(new_n892_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n616_), .A3(new_n892_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n892_), .A2(new_n616_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n309_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n907_), .A2(new_n326_), .B1(new_n891_), .B2(new_n909_), .ZN(G1350gat));
  NAND2_X1  g709(.A1(new_n893_), .A2(new_n586_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(G190gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n893_), .A2(new_n310_), .A3(new_n614_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1351gat));
  NAND4_X1  g713(.A1(new_n425_), .A2(new_n257_), .A3(new_n301_), .A4(new_n622_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n831_), .B2(new_n841_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n467_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(KEYINPUT126), .B2(new_n281_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT126), .B(G197gat), .Z(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n917_), .B2(new_n919_), .ZN(G1352gat));
  AND2_X1   g719(.A1(new_n916_), .A2(new_n720_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(G204gat), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n273_), .B2(new_n921_), .ZN(G1353gat));
  AOI21_X1  g722(.A(new_n600_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n916_), .A2(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n925_), .B(new_n926_), .Z(G1354gat));
  NOR2_X1   g726(.A1(new_n837_), .A2(G218gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n916_), .A2(new_n928_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n916_), .A2(new_n586_), .ZN(new_n930_));
  INV_X1    g729(.A(G218gat), .ZN(new_n931_));
  OAI211_X1 g730(.A(KEYINPUT127), .B(new_n929_), .C1(new_n930_), .C2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933_));
  INV_X1    g732(.A(new_n929_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n931_), .B1(new_n916_), .B2(new_n586_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n933_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n932_), .A2(new_n936_), .ZN(G1355gat));
endmodule


