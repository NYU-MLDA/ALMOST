//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT70), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n202_), .B(KEYINPUT70), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT11), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT69), .B(G71gat), .ZN(new_n208_));
  INV_X1    g007(.A(G78gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n205_), .A2(new_n207_), .A3(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n207_), .A2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G231gat), .A2(G233gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT77), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217_));
  INV_X1    g016(.A(G1gat), .ZN(new_n218_));
  INV_X1    g017(.A(G8gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT14), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G1gat), .B(G8gat), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n221_), .B(new_n222_), .Z(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n216_), .B(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G127gat), .B(G155gat), .Z(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT16), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G183gat), .B(G211gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n225_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT78), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(KEYINPUT78), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n229_), .B(new_n230_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n225_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT37), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G29gat), .B(G36gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT74), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT15), .ZN(new_n245_));
  AOI211_X1 g044(.A(G99gat), .B(G106gat), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(KEYINPUT67), .B2(KEYINPUT7), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT66), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G99gat), .A2(G106gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT6), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G85gat), .B(G92gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n253_), .A2(KEYINPUT68), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT8), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT65), .B(G85gat), .ZN(new_n257_));
  INV_X1    g056(.A(G92gat), .ZN(new_n258_));
  OR3_X1    g057(.A1(new_n257_), .A2(KEYINPUT9), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n253_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT9), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT10), .B(G99gat), .Z(new_n262_));
  INV_X1    g061(.A(G106gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n259_), .A2(new_n261_), .A3(new_n264_), .A4(new_n251_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n256_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n245_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n256_), .A2(new_n244_), .A3(new_n265_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G232gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT34), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n267_), .B(new_n268_), .C1(KEYINPUT35), .C2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(KEYINPUT35), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n271_), .B(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT76), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT36), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G190gat), .B(G218gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT75), .ZN(new_n278_));
  XOR2_X1   g077(.A(G134gat), .B(G162gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n275_), .A2(new_n276_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  OAI22_X1  g081(.A1(new_n274_), .A2(KEYINPUT76), .B1(KEYINPUT36), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n274_), .A2(KEYINPUT36), .A3(new_n282_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n240_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n284_), .A2(new_n240_), .A3(new_n285_), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n239_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G230gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT64), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n213_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n266_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n266_), .A2(new_n292_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n293_), .B1(new_n295_), .B2(KEYINPUT12), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT12), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n298_), .A2(KEYINPUT71), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(KEYINPUT71), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n291_), .B(new_n296_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT72), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n290_), .B1(new_n295_), .B2(new_n293_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n298_), .B(KEYINPUT71), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n291_), .A4(new_n296_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G120gat), .B(G148gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT5), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G176gat), .B(G204gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n302_), .A2(new_n306_), .A3(new_n303_), .A4(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT13), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(KEYINPUT13), .A3(new_n314_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(KEYINPUT73), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n318_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n288_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT79), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n326_));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT84), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n327_), .B(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n332_), .B2(new_n329_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OR3_X1    g133(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n336_), .B(KEYINPUT83), .Z(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT25), .B(G183gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT82), .ZN(new_n342_));
  INV_X1    g141(.A(G190gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT26), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n343_), .A2(KEYINPUT26), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n341_), .B(new_n344_), .C1(new_n345_), .C2(new_n342_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n334_), .A2(new_n335_), .A3(new_n340_), .A4(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n328_), .A2(KEYINPUT23), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n332_), .B2(KEYINPUT23), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT22), .B(G169gat), .ZN(new_n353_));
  INV_X1    g152(.A(G176gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n337_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G43gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n347_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n347_), .B2(new_n357_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n326_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n347_), .A2(new_n357_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n359_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n326_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n360_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G127gat), .B(G134gat), .Z(new_n369_));
  XOR2_X1   g168(.A(G113gat), .B(G120gat), .Z(new_n370_));
  XOR2_X1   g169(.A(new_n369_), .B(new_n370_), .Z(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(G15gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT30), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n371_), .B(new_n375_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n363_), .A2(new_n368_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n363_), .B2(new_n368_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G211gat), .B(G218gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G197gat), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n383_), .A2(KEYINPUT89), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(KEYINPUT89), .ZN(new_n385_));
  INV_X1    g184(.A(G204gat), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT90), .B(G204gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(G197gat), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT21), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n382_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT91), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n388_), .B2(G197gat), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(G204gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n386_), .A2(KEYINPUT90), .ZN(new_n396_));
  OAI211_X1 g195(.A(KEYINPUT91), .B(new_n383_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n386_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT92), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT21), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n399_), .B2(KEYINPUT21), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n391_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  OR3_X1    g202(.A1(new_n389_), .A2(new_n390_), .A3(new_n381_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OR2_X1    g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT3), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT2), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n407_), .B2(KEYINPUT1), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT1), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n417_), .A2(KEYINPUT86), .A3(G155gat), .A4(G162gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n407_), .A2(KEYINPUT1), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n416_), .A2(new_n418_), .A3(new_n419_), .A4(new_n406_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G141gat), .B(G148gat), .Z(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(KEYINPUT87), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT87), .B1(new_n420_), .B2(new_n421_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n414_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n405_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G228gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n420_), .A2(new_n421_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n413_), .B1(new_n434_), .B2(new_n422_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT29), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT88), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n425_), .A2(new_n438_), .A3(KEYINPUT29), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n428_), .A2(new_n430_), .B1(new_n431_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT94), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n443_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n435_), .A2(new_n436_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G22gat), .B(G50gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT28), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n448_), .B(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .A4(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n447_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n446_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n451_), .ZN(new_n455_));
  OAI22_X1  g254(.A1(new_n453_), .A2(new_n444_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G225gat), .A2(G233gat), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n459_), .B(KEYINPUT96), .Z(new_n460_));
  NAND2_X1  g259(.A1(new_n425_), .A2(new_n371_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n371_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n435_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n460_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n461_), .A2(new_n463_), .A3(KEYINPUT4), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT97), .B(KEYINPUT4), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n425_), .A2(new_n371_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT98), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT98), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n425_), .A2(new_n469_), .A3(new_n371_), .A4(new_n466_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n464_), .B1(new_n471_), .B2(new_n460_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G1gat), .B(G29gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G85gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT0), .B(G57gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OR3_X1    g276(.A1(new_n472_), .A2(KEYINPUT33), .A3(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT33), .B1(new_n472_), .B2(new_n477_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n334_), .A2(new_n351_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n336_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n335_), .B1(new_n482_), .B2(new_n338_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT26), .B(G190gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n341_), .B2(new_n484_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n481_), .A2(new_n356_), .B1(new_n349_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n405_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n403_), .A2(new_n404_), .A3(new_n357_), .A4(new_n347_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT20), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G226gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT19), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT95), .Z(new_n493_));
  NAND3_X1  g292(.A1(new_n403_), .A2(new_n404_), .A3(new_n486_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n494_), .A2(KEYINPUT20), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n492_), .B1(new_n405_), .B2(new_n364_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n490_), .A2(new_n493_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G8gat), .B(G36gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT18), .ZN(new_n499_));
  XOR2_X1   g298(.A(G64gat), .B(G92gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n497_), .A2(new_n501_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n461_), .A2(new_n463_), .A3(new_n460_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n477_), .B(new_n504_), .C1(new_n471_), .C2(new_n460_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n480_), .A2(new_n502_), .A3(new_n503_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(KEYINPUT32), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n497_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n472_), .A2(new_n477_), .ZN(new_n509_));
  AOI211_X1 g308(.A(new_n476_), .B(new_n464_), .C1(new_n471_), .C2(new_n460_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n493_), .ZN(new_n512_));
  AND4_X1   g311(.A1(KEYINPUT20), .A2(new_n488_), .A3(new_n512_), .A4(new_n489_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n494_), .A2(KEYINPUT20), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT99), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n494_), .A2(KEYINPUT99), .A3(KEYINPUT20), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n405_), .A2(new_n364_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n513_), .B1(new_n519_), .B2(new_n492_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT100), .B1(new_n520_), .B2(new_n507_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT100), .ZN(new_n522_));
  INV_X1    g321(.A(new_n507_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n492_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n514_), .A2(new_n515_), .B1(new_n405_), .B2(new_n364_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n524_), .B1(new_n525_), .B2(new_n517_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n522_), .B(new_n523_), .C1(new_n526_), .C2(new_n513_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n511_), .B1(new_n521_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n506_), .B1(new_n528_), .B2(KEYINPUT101), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT101), .ZN(new_n530_));
  AOI211_X1 g329(.A(new_n530_), .B(new_n511_), .C1(new_n521_), .C2(new_n527_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n458_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n503_), .A2(new_n502_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT27), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n536_), .B(KEYINPUT102), .C1(new_n501_), .C2(new_n520_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n509_), .A2(new_n510_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT102), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n520_), .A2(new_n501_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n536_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n538_), .A2(new_n539_), .A3(new_n457_), .A4(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n380_), .B1(new_n532_), .B2(new_n544_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n509_), .A2(new_n379_), .A3(new_n510_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n546_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n547_), .A2(new_n543_), .A3(new_n535_), .A4(new_n537_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT103), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n244_), .B(new_n223_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT80), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n245_), .A2(new_n224_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n244_), .A2(new_n223_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n552_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G113gat), .B(G141gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT81), .ZN(new_n561_));
  XOR2_X1   g360(.A(G169gat), .B(G197gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n550_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n325_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n539_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n218_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT38), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n284_), .A2(new_n285_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n550_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n322_), .A2(new_n319_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n567_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n239_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(G1gat), .B1(new_n581_), .B2(new_n539_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n572_), .A2(new_n573_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n574_), .A2(new_n582_), .A3(new_n583_), .ZN(G1324gat));
  XNOR2_X1  g383(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n538_), .A2(new_n543_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G8gat), .B1(new_n581_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT104), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(KEYINPUT104), .B(G8gat), .C1(new_n581_), .C2(new_n588_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(KEYINPUT39), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n587_), .A2(new_n219_), .ZN(new_n595_));
  OAI22_X1  g394(.A1(new_n591_), .A2(KEYINPUT39), .B1(new_n569_), .B2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n586_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n569_), .A2(new_n595_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n589_), .A2(new_n590_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n593_), .A3(new_n585_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n602_), .ZN(G1325gat));
  OAI21_X1  g402(.A(G15gat), .B1(new_n581_), .B2(new_n379_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT41), .Z(new_n605_));
  NAND3_X1  g404(.A1(new_n570_), .A2(new_n373_), .A3(new_n380_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(G1326gat));
  XNOR2_X1  g406(.A(new_n457_), .B(KEYINPUT106), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G22gat), .B1(new_n581_), .B2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT42), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n609_), .A2(G22gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n611_), .B1(new_n569_), .B2(new_n612_), .ZN(G1327gat));
  INV_X1    g412(.A(new_n578_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n237_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(new_n576_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n568_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(G29gat), .B1(new_n618_), .B2(new_n571_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n286_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n284_), .A2(new_n240_), .A3(new_n285_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT43), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n622_), .B(new_n625_), .C1(new_n545_), .C2(new_n549_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n578_), .A2(new_n579_), .A3(new_n615_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(KEYINPUT44), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT44), .B1(new_n627_), .B2(new_n628_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n571_), .A2(G29gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n619_), .B1(new_n631_), .B2(new_n632_), .ZN(G1328gat));
  INV_X1    g432(.A(G36gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n587_), .A2(new_n634_), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n617_), .A2(KEYINPUT45), .A3(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT45), .B1(new_n617_), .B2(new_n635_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n629_), .A2(new_n630_), .A3(new_n588_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n634_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n638_), .B(KEYINPUT46), .C1(new_n639_), .C2(new_n634_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1329gat));
  AOI21_X1  g443(.A(G43gat), .B1(new_n618_), .B2(new_n380_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n380_), .A2(G43gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n631_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT47), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1330gat));
  AOI21_X1  g448(.A(G50gat), .B1(new_n618_), .B2(new_n608_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n457_), .A2(G50gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n631_), .B2(new_n651_), .ZN(G1331gat));
  NAND2_X1  g451(.A1(new_n550_), .A2(new_n579_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n550_), .A2(KEYINPUT107), .A3(new_n579_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(new_n578_), .A3(new_n288_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G57gat), .B1(new_n658_), .B2(new_n571_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n614_), .A2(new_n567_), .A3(new_n239_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(KEYINPUT108), .B(G57gat), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n660_), .A2(new_n571_), .A3(new_n577_), .A4(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT109), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n659_), .A2(new_n663_), .ZN(G1332gat));
  NAND2_X1  g463(.A1(new_n660_), .A2(new_n577_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G64gat), .B1(new_n665_), .B2(new_n588_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT48), .ZN(new_n667_));
  INV_X1    g466(.A(G64gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n658_), .A2(new_n668_), .A3(new_n587_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1333gat));
  OAI21_X1  g469(.A(G71gat), .B1(new_n665_), .B2(new_n379_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT49), .ZN(new_n672_));
  INV_X1    g471(.A(G71gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n658_), .A2(new_n673_), .A3(new_n380_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1334gat));
  OAI21_X1  g474(.A(G78gat), .B1(new_n665_), .B2(new_n609_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT50), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n658_), .A2(new_n209_), .A3(new_n608_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1335gat));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n578_), .A2(new_n616_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n680_), .B1(new_n657_), .B2(new_n682_), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT110), .B(new_n681_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n571_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(G85gat), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n624_), .A2(KEYINPUT111), .A3(new_n626_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT111), .B1(new_n624_), .B2(new_n626_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n239_), .A2(new_n579_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n689_), .A2(new_n614_), .A3(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n539_), .A2(new_n257_), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n685_), .A2(new_n686_), .B1(new_n691_), .B2(new_n692_), .ZN(G1336gat));
  NAND2_X1  g492(.A1(new_n657_), .A2(new_n682_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT110), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n657_), .A2(new_n680_), .A3(new_n682_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n588_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT112), .B1(new_n697_), .B2(G92gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n587_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT112), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n258_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n588_), .A2(new_n258_), .ZN(new_n702_));
  AOI22_X1  g501(.A1(new_n698_), .A2(new_n701_), .B1(new_n691_), .B2(new_n702_), .ZN(G1337gat));
  AND2_X1   g502(.A1(new_n380_), .A2(new_n262_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n614_), .A2(new_n690_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n380_), .B(new_n706_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT113), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(G99gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n707_), .B2(G99gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT51), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n713_), .B(new_n705_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1338gat));
  NOR2_X1   g514(.A1(new_n458_), .A2(G106gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n690_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n578_), .A2(new_n457_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT114), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n627_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G106gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n720_), .B2(new_n627_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n723_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n725_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n719_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n263_), .B1(new_n728_), .B2(new_n721_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n724_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n717_), .B1(new_n726_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n717_), .B(new_n733_), .C1(new_n726_), .C2(new_n731_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1339gat));
  NAND3_X1  g536(.A1(new_n556_), .A2(new_n557_), .A3(new_n553_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n564_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n559_), .A2(new_n564_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n314_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n302_), .A2(new_n742_), .A3(new_n306_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n304_), .A2(new_n296_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n290_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n745_), .B1(new_n742_), .B2(new_n301_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n311_), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n302_), .A2(new_n742_), .A3(new_n306_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(new_n745_), .C1(new_n742_), .C2(new_n301_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT56), .B1(new_n751_), .B2(new_n311_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n741_), .B1(new_n749_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT58), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT58), .B(new_n741_), .C1(new_n749_), .C2(new_n752_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n622_), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n567_), .A2(new_n314_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n747_), .A2(new_n748_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n311_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n315_), .A2(new_n740_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n576_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT57), .B(new_n576_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n757_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n239_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n287_), .A2(new_n286_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(new_n579_), .A3(new_n615_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(new_n320_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n320_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n769_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n288_), .A2(new_n579_), .A3(new_n773_), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n768_), .A2(new_n777_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n587_), .A2(new_n539_), .A3(new_n379_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n458_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n776_), .B1(new_n767_), .B2(new_n239_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(new_n457_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(KEYINPUT59), .A3(new_n779_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(G113gat), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n579_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  INV_X1    g588(.A(new_n779_), .ZN(new_n790_));
  NOR4_X1   g589(.A1(new_n783_), .A2(new_n457_), .A3(new_n579_), .A4(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n791_), .B2(G113gat), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT118), .B(new_n787_), .C1(new_n780_), .C2(new_n579_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n786_), .A2(new_n788_), .B1(new_n792_), .B2(new_n793_), .ZN(G1340gat));
  INV_X1    g593(.A(new_n780_), .ZN(new_n795_));
  INV_X1    g594(.A(G120gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n614_), .B2(KEYINPUT60), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n795_), .B(new_n797_), .C1(KEYINPUT60), .C2(new_n796_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n614_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n796_), .ZN(G1341gat));
  INV_X1    g599(.A(G127gat), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n239_), .A2(new_n801_), .ZN(new_n802_));
  NOR4_X1   g601(.A1(new_n783_), .A2(new_n457_), .A3(new_n239_), .A4(new_n790_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT119), .B1(new_n803_), .B2(G127gat), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n801_), .C1(new_n780_), .C2(new_n239_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n786_), .A2(new_n802_), .B1(new_n804_), .B2(new_n806_), .ZN(G1342gat));
  INV_X1    g606(.A(G134gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n795_), .A2(new_n808_), .A3(new_n575_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n770_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n808_), .ZN(G1343gat));
  NAND3_X1  g610(.A1(new_n457_), .A2(new_n571_), .A3(new_n379_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n783_), .A2(new_n587_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n567_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n578_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT120), .B(G148gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1345gat));
  NAND2_X1  g617(.A1(new_n813_), .A2(new_n615_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT61), .B(G155gat), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1346gat));
  INV_X1    g620(.A(G162gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n813_), .A2(new_n822_), .A3(new_n575_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n813_), .A2(new_n622_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n822_), .ZN(G1347gat));
  NAND2_X1  g624(.A1(new_n587_), .A2(new_n546_), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT121), .Z(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n783_), .A2(new_n608_), .A3(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(new_n353_), .A3(new_n567_), .ZN(new_n830_));
  INV_X1    g629(.A(G169gat), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n783_), .A2(new_n608_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n827_), .A2(new_n567_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT122), .Z(new_n834_));
  AOI21_X1  g633(.A(new_n831_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n835_), .A2(new_n836_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n837_), .B2(new_n838_), .ZN(G1348gat));
  NAND3_X1  g638(.A1(new_n829_), .A2(new_n354_), .A3(new_n578_), .ZN(new_n840_));
  NOR4_X1   g639(.A1(new_n783_), .A2(new_n457_), .A3(new_n614_), .A4(new_n828_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n354_), .B2(new_n841_), .ZN(G1349gat));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n843_));
  INV_X1    g642(.A(new_n341_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n828_), .A2(new_n239_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n832_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G183gat), .B1(new_n784_), .B2(new_n845_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n843_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n784_), .A2(new_n845_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT123), .B(new_n846_), .C1(new_n850_), .C2(G183gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1350gat));
  NAND2_X1  g651(.A1(new_n575_), .A2(new_n484_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT125), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n829_), .A2(new_n854_), .ZN(new_n855_));
  AOI211_X1 g654(.A(KEYINPUT124), .B(new_n343_), .C1(new_n829_), .C2(new_n622_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n832_), .A2(new_n622_), .A3(new_n827_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(G190gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n856_), .B2(new_n859_), .ZN(G1351gat));
  NOR4_X1   g659(.A1(new_n588_), .A2(new_n571_), .A3(new_n458_), .A4(new_n380_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n778_), .A2(KEYINPUT126), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT126), .ZN(new_n863_));
  INV_X1    g662(.A(new_n861_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n783_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n579_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(new_n383_), .ZN(G1352gat));
  NAND2_X1  g666(.A1(new_n862_), .A2(new_n865_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G204gat), .B1(new_n868_), .B2(new_n578_), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n388_), .B(new_n614_), .C1(new_n862_), .C2(new_n865_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1353gat));
  AOI21_X1  g670(.A(new_n239_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT127), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n873_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n868_), .A2(new_n872_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n872_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n878_), .B(new_n875_), .C1(new_n862_), .C2(new_n865_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1354gat));
  INV_X1    g679(.A(G218gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n868_), .A2(new_n881_), .A3(new_n575_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n770_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(new_n883_), .ZN(G1355gat));
endmodule


