//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n945_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT72), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT34), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT35), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(KEYINPUT6), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(KEYINPUT66), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n212_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(KEYINPUT66), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(KEYINPUT6), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(G99gat), .A4(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT7), .ZN(new_n222_));
  INV_X1    g021(.A(G99gat), .ZN(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n211_), .B1(new_n221_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT8), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n225_), .A2(KEYINPUT67), .A3(new_n226_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(KEYINPUT8), .B(new_n211_), .C1(new_n234_), .C2(new_n221_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n221_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT10), .B(G99gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT64), .B(G106gat), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT9), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n208_), .A2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n240_), .B(new_n242_), .C1(new_n211_), .C2(new_n241_), .ZN(new_n243_));
  OR2_X1    g042(.A1(G85gat), .A2(G92gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n241_), .B1(new_n244_), .B2(new_n208_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n242_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT65), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n236_), .A2(new_n239_), .A3(new_n243_), .A4(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n230_), .A2(new_n235_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G50gat), .ZN(new_n250_));
  OR2_X1    g049(.A1(G29gat), .A2(G36gat), .ZN(new_n251_));
  INV_X1    g050(.A(G43gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G29gat), .A2(G36gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n252_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n250_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n251_), .A2(new_n253_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G43gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(G50gat), .A3(new_n254_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n257_), .A2(KEYINPUT15), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT15), .B1(new_n257_), .B2(new_n260_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n249_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n205_), .A2(new_n206_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n260_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n249_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n263_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n239_), .A2(new_n220_), .A3(new_n217_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n247_), .A2(new_n243_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n269_), .A2(new_n270_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n255_), .A2(new_n250_), .A3(new_n256_), .ZN(new_n272_));
  AOI21_X1  g071(.A(G50gat), .B1(new_n259_), .B2(new_n254_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n271_), .A2(new_n235_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT73), .B1(new_n275_), .B2(new_n264_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n202_), .B(new_n207_), .C1(new_n268_), .C2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n266_), .A2(new_n267_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(KEYINPUT73), .A3(new_n264_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n263_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n202_), .B1(new_n281_), .B2(new_n207_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT36), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT75), .B(G134gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G162gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G190gat), .B(G218gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  INV_X1    g087(.A(new_n207_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n263_), .A2(new_n275_), .A3(new_n289_), .A4(new_n264_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n283_), .A2(new_n284_), .A3(new_n288_), .A4(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n207_), .B1(new_n268_), .B2(new_n276_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT74), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n277_), .A3(new_n290_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n288_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT36), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(KEYINPUT36), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT37), .B1(new_n291_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n291_), .A2(new_n299_), .A3(KEYINPUT37), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G127gat), .B(G155gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(G183gat), .B(G211gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT17), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT77), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G15gat), .B(G22gat), .ZN(new_n311_));
  INV_X1    g110(.A(G1gat), .ZN(new_n312_));
  INV_X1    g111(.A(G8gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT14), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G1gat), .B(G8gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G231gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G57gat), .ZN(new_n320_));
  INV_X1    g119(.A(G64gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G57gat), .A2(G64gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT11), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G71gat), .B(G78gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT11), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n322_), .A2(new_n328_), .A3(new_n323_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n326_), .A3(KEYINPUT11), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n319_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n310_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n330_), .A2(KEYINPUT68), .A3(new_n331_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n319_), .B(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n308_), .A2(KEYINPUT17), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n309_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n335_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n303_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT78), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n330_), .A2(KEYINPUT68), .A3(new_n331_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT68), .B1(new_n330_), .B2(new_n331_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n249_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT12), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n249_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n339_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G230gat), .A2(G233gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n249_), .A2(KEYINPUT12), .A3(new_n333_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT69), .B1(new_n249_), .B2(new_n348_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n271_), .A2(new_n339_), .A3(new_n359_), .A4(new_n235_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n349_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n354_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(KEYINPUT70), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT70), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n358_), .A2(new_n360_), .B1(new_n348_), .B2(new_n249_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n365_), .B1(new_n366_), .B2(new_n354_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n357_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G120gat), .B(G148gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(G204gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT5), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G176gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  AOI211_X1 g173(.A(new_n372_), .B(new_n357_), .C1(new_n364_), .C2(new_n367_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT13), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n376_), .B1(KEYINPUT71), .B2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT79), .B1(new_n265_), .B2(new_n317_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n265_), .A2(new_n317_), .A3(KEYINPUT79), .ZN(new_n384_));
  INV_X1    g183(.A(new_n317_), .ZN(new_n385_));
  OAI22_X1  g184(.A1(new_n383_), .A2(new_n384_), .B1(new_n385_), .B2(new_n274_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G229gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  OR3_X1    g188(.A1(new_n265_), .A2(new_n317_), .A3(KEYINPUT79), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n382_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n317_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT80), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n394_), .B(new_n317_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n391_), .A2(new_n393_), .A3(new_n387_), .A4(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G113gat), .B(G141gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G197gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT81), .ZN(new_n399_));
  INV_X1    g198(.A(G169gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n389_), .A2(new_n396_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n389_), .B2(new_n396_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n381_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G211gat), .B(G218gat), .ZN(new_n409_));
  INV_X1    g208(.A(G197gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT91), .B1(new_n410_), .B2(G204gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(KEYINPUT21), .A3(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G197gat), .B(G204gat), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n409_), .A2(KEYINPUT21), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n413_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G183gat), .A2(G190gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT23), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT24), .ZN(new_n423_));
  INV_X1    g222(.A(G176gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n400_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n422_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G190gat), .ZN(new_n428_));
  INV_X1    g227(.A(G183gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT25), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT82), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT25), .B(G183gat), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n428_), .B(new_n432_), .C1(new_n433_), .C2(new_n431_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n425_), .A2(KEYINPUT24), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n427_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n420_), .B(new_n421_), .C1(G183gat), .C2(G190gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT22), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n439_), .B(G169gat), .C1(new_n440_), .C2(KEYINPUT83), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT22), .B1(new_n400_), .B2(KEYINPUT84), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n424_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n426_), .A2(KEYINPUT83), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n438_), .A2(new_n443_), .A3(new_n444_), .A4(new_n435_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n417_), .A2(new_n437_), .A3(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT22), .B(G169gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n424_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n438_), .A3(new_n435_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n422_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n423_), .A2(KEYINPUT95), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT24), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n426_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n425_), .A2(new_n452_), .A3(new_n454_), .A4(new_n435_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G183gat), .ZN(new_n459_));
  AND2_X1   g258(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n430_), .B(new_n459_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT96), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n457_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n463_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n451_), .B(new_n456_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT97), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n457_), .A2(new_n462_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT96), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n457_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT97), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n451_), .A4(new_n456_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n450_), .B1(new_n467_), .B2(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(KEYINPUT20), .B(new_n446_), .C1(new_n474_), .C2(new_n417_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT94), .ZN(new_n477_));
  AND2_X1   g276(.A1(G226gat), .A2(G233gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n475_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n422_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n472_), .B1(new_n482_), .B2(new_n456_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n466_), .A2(KEYINPUT97), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n417_), .B(new_n449_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT98), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT20), .ZN(new_n487_));
  INV_X1    g286(.A(new_n417_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n437_), .A2(new_n445_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT98), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n474_), .A2(new_n491_), .A3(new_n417_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n486_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n481_), .B1(new_n480_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT18), .B(G64gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G92gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G8gat), .B(G36gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n496_), .B(new_n497_), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT32), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n449_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n488_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n502_), .A2(KEYINPUT20), .A3(new_n480_), .A4(new_n446_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n466_), .A2(new_n417_), .A3(new_n449_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n490_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n479_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n499_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT103), .ZN(new_n508_));
  OAI22_X1  g307(.A1(new_n494_), .A2(new_n500_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n493_), .A2(new_n480_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n481_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(KEYINPUT103), .A3(new_n499_), .ZN(new_n513_));
  INV_X1    g312(.A(G141gat), .ZN(new_n514_));
  INV_X1    g313(.A(G148gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G141gat), .A2(G148gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G155gat), .A2(G162gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT1), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520_));
  INV_X1    g319(.A(G155gat), .ZN(new_n521_));
  INV_X1    g320(.A(G162gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n516_), .B(new_n517_), .C1(new_n519_), .C2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n527_));
  NOR2_X1   g326(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(new_n528_), .B2(new_n517_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT3), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(KEYINPUT88), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n529_), .A2(new_n530_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n523_), .A2(new_n524_), .A3(new_n518_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n534_), .A2(KEYINPUT89), .A3(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT89), .B1(new_n534_), .B2(new_n535_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n526_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G127gat), .B(G134gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G113gat), .ZN(new_n540_));
  OR2_X1    g339(.A1(G127gat), .A2(G134gat), .ZN(new_n541_));
  INV_X1    g340(.A(G113gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G127gat), .A2(G134gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n540_), .A2(G120gat), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(G120gat), .B1(new_n540_), .B2(new_n544_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n538_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n547_), .B(new_n526_), .C1(new_n537_), .C2(new_n536_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(KEYINPUT99), .A3(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n536_), .A2(new_n537_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT99), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n526_), .A4(new_n547_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n554_), .A3(KEYINPUT4), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT4), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n549_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G225gat), .A2(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n551_), .A2(new_n554_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n559_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT0), .B(G57gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(G85gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(G1gat), .B(G29gat), .Z(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n561_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n563_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n559_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n567_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n509_), .A2(new_n513_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n512_), .A2(new_n498_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT101), .B(KEYINPUT33), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n569_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n498_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n494_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n568_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT102), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n562_), .B(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n580_), .B1(new_n582_), .B2(new_n559_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n575_), .A2(new_n577_), .A3(new_n579_), .A4(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT33), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n585_), .B1(new_n569_), .B2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n570_), .A2(new_n571_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n588_), .A2(KEYINPUT100), .A3(KEYINPUT33), .A4(new_n568_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n574_), .B1(new_n584_), .B2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G78gat), .B(G106gat), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n417_), .B1(new_n538_), .B2(KEYINPUT29), .ZN(new_n594_));
  INV_X1    g393(.A(G228gat), .ZN(new_n595_));
  INV_X1    g394(.A(G233gat), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  AOI211_X1 g398(.A(new_n597_), .B(new_n417_), .C1(new_n538_), .C2(KEYINPUT29), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n593_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT92), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n538_), .A2(KEYINPUT29), .ZN(new_n603_));
  XOR2_X1   g402(.A(G22gat), .B(G50gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n603_), .B(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n594_), .A2(new_n598_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n600_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n592_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n602_), .A2(new_n607_), .B1(new_n610_), .B2(new_n601_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n610_), .A2(new_n607_), .A3(new_n601_), .A4(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT86), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT30), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n437_), .A2(new_n445_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n618_), .B1(new_n437_), .B2(new_n445_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n548_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n489_), .A2(KEYINPUT30), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n547_), .A3(new_n619_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G71gat), .B(G99gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G227gat), .A2(G233gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n622_), .A2(new_n624_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n628_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G15gat), .B(G43gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n630_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n622_), .A2(new_n624_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n627_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n634_), .B1(new_n638_), .B2(new_n629_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n617_), .B1(new_n636_), .B2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n635_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n634_), .A3(new_n629_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(KEYINPUT86), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n616_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT27), .B1(new_n575_), .B2(new_n579_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n578_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT27), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n498_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n646_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n640_), .B(new_n643_), .C1(new_n611_), .C2(new_n614_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n602_), .A2(new_n607_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n610_), .A2(new_n601_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n641_), .A2(new_n642_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n613_), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n573_), .B1(new_n652_), .B2(new_n657_), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n591_), .A2(new_n645_), .B1(new_n651_), .B2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n408_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n345_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n312_), .A3(new_n573_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT38), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n291_), .A2(new_n299_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n343_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n660_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n573_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G1gat), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n663_), .A2(new_n670_), .ZN(G1324gat));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672_));
  INV_X1    g471(.A(new_n651_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n660_), .A2(new_n667_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(G8gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n675_), .B1(new_n674_), .B2(G8gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n672_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n678_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(KEYINPUT105), .A3(new_n676_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n681_), .A3(KEYINPUT39), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n661_), .A2(new_n313_), .A3(new_n673_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n672_), .B(new_n684_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n683_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1325gat));
  INV_X1    g487(.A(new_n644_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G15gat), .B1(new_n668_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT41), .Z(new_n691_));
  INV_X1    g490(.A(G15gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n661_), .A2(new_n692_), .A3(new_n644_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1326gat));
  OAI21_X1  g493(.A(G22gat), .B1(new_n668_), .B2(new_n615_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT42), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n615_), .A2(G22gat), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT106), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n661_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1327gat));
  NOR2_X1   g499(.A1(new_n659_), .A2(new_n664_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n381_), .A2(new_n343_), .A3(new_n407_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n573_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n591_), .A2(new_n645_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n651_), .A2(new_n658_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n303_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n291_), .A2(KEYINPUT37), .A3(new_n299_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(new_n300_), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT43), .B1(new_n659_), .B2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n702_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(KEYINPUT44), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(KEYINPUT44), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n715_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n669_), .B(new_n716_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n706_), .B1(new_n721_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g521(.A(G36gat), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n701_), .A2(new_n703_), .A3(new_n723_), .A4(new_n673_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT45), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n673_), .B1(new_n715_), .B2(KEYINPUT44), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n725_), .B1(new_n727_), .B2(new_n723_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT108), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(KEYINPUT46), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n728_), .B2(KEYINPUT109), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT109), .B1(new_n728_), .B2(KEYINPUT108), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n733_), .B2(new_n734_), .ZN(G1329gat));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n719_), .A2(new_n720_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n716_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n656_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(new_n252_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n252_), .B1(new_n704_), .B2(new_n689_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n736_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n741_), .A2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT110), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(KEYINPUT47), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n750_), .ZN(G1330gat));
  NAND3_X1  g550(.A1(new_n737_), .A2(new_n616_), .A3(new_n738_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n752_), .A2(KEYINPUT111), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(KEYINPUT111), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(G50gat), .A3(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n705_), .A2(new_n250_), .A3(new_n616_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1331gat));
  NOR2_X1   g556(.A1(new_n381_), .A2(new_n407_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n759_), .A2(new_n666_), .A3(new_n659_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n761_), .A2(new_n320_), .A3(new_n669_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n345_), .A2(new_n709_), .A3(new_n758_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n573_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n764_), .B2(new_n320_), .ZN(G1332gat));
  AOI21_X1  g564(.A(new_n321_), .B1(new_n760_), .B2(new_n673_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT48), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(new_n321_), .A3(new_n673_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1333gat));
  INV_X1    g568(.A(G71gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n760_), .B2(new_n644_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT49), .Z(new_n772_));
  NAND3_X1  g571(.A1(new_n763_), .A2(new_n770_), .A3(new_n644_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1334gat));
  OAI21_X1  g573(.A(G78gat), .B1(new_n761_), .B2(new_n615_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT50), .ZN(new_n776_));
  INV_X1    g575(.A(G78gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n763_), .A2(new_n777_), .A3(new_n616_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT112), .ZN(G1335gat));
  NOR3_X1   g579(.A1(new_n381_), .A2(new_n665_), .A3(new_n407_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n701_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n573_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n710_), .B1(new_n709_), .B2(new_n303_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n659_), .A2(KEYINPUT43), .A3(new_n713_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n781_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT113), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n758_), .A2(new_n343_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n789_), .A2(new_n794_), .A3(new_n669_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n784_), .B1(new_n795_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g595(.A(G92gat), .B1(new_n783_), .B2(new_n673_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n789_), .A2(new_n794_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n673_), .A2(G92gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n798_), .B2(new_n799_), .ZN(G1337gat));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT51), .ZN(new_n802_));
  OR3_X1    g601(.A1(new_n782_), .A2(new_n237_), .A3(new_n739_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n788_), .A2(new_n644_), .A3(new_n793_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n804_), .A2(new_n805_), .A3(G99gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n804_), .B2(G99gat), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n802_), .B(new_n803_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n801_), .A2(KEYINPUT51), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n804_), .A2(G99gat), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT114), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n804_), .A2(new_n805_), .A3(G99gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n809_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n810_), .A2(new_n816_), .ZN(G1338gat));
  OR3_X1    g616(.A1(new_n782_), .A2(new_n238_), .A3(new_n615_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n791_), .A2(new_n616_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(G106gat), .ZN(new_n821_));
  AOI211_X1 g620(.A(KEYINPUT52), .B(new_n224_), .C1(new_n791_), .C2(new_n616_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n344_), .A2(new_n825_), .A3(new_n406_), .A4(new_n381_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n713_), .A2(new_n665_), .A3(new_n406_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n381_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT54), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n826_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n386_), .A2(new_n387_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n391_), .A2(new_n393_), .A3(new_n388_), .A4(new_n395_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n401_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n403_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n403_), .A2(new_n833_), .A3(KEYINPUT116), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT117), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n375_), .A2(new_n406_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n357_), .A2(KEYINPUT55), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n361_), .A2(new_n351_), .A3(new_n355_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n363_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n356_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n842_), .A2(new_n844_), .A3(new_n846_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n847_), .A2(KEYINPUT56), .A3(new_n372_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT56), .B1(new_n847_), .B2(new_n372_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n841_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n838_), .B(new_n851_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n840_), .A2(new_n850_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n664_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n375_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(new_n838_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n859_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n303_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n853_), .A2(KEYINPUT57), .A3(new_n664_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n856_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n864_), .A2(KEYINPUT118), .A3(new_n343_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT118), .B1(new_n864_), .B2(new_n343_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n830_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n673_), .A2(new_n669_), .A3(new_n657_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n864_), .A2(new_n343_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n830_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n869_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT59), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n870_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(G113gat), .A3(new_n407_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n542_), .B1(new_n873_), .B2(new_n406_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1340gat));
  NAND3_X1  g677(.A1(new_n870_), .A2(new_n828_), .A3(new_n874_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT119), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n870_), .A2(new_n881_), .A3(new_n828_), .A4(new_n874_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(G120gat), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n873_), .ZN(new_n884_));
  INV_X1    g683(.A(G120gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n381_), .B2(KEYINPUT60), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n884_), .B(new_n886_), .C1(KEYINPUT60), .C2(new_n885_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n887_), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n343_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n870_), .A2(new_n874_), .A3(new_n890_), .ZN(new_n891_));
  OAI211_X1 g690(.A(KEYINPUT120), .B(new_n889_), .C1(new_n873_), .C2(new_n343_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n889_), .B1(new_n873_), .B2(new_n343_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n892_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT121), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n891_), .A2(new_n898_), .A3(new_n895_), .A4(new_n892_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1342gat));
  INV_X1    g699(.A(new_n664_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G134gat), .B1(new_n884_), .B2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n303_), .A2(G134gat), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT122), .Z(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n875_), .B2(new_n904_), .ZN(G1343gat));
  AOI21_X1  g704(.A(new_n652_), .B1(new_n871_), .B2(new_n830_), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n906_), .A2(new_n573_), .A3(new_n651_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n407_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n828_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT123), .B(G148gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1345gat));
  NAND2_X1  g711(.A1(new_n907_), .A2(new_n665_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT61), .B(G155gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1346gat));
  AOI21_X1  g714(.A(G162gat), .B1(new_n907_), .B2(new_n901_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n713_), .A2(new_n522_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n907_), .B2(new_n917_), .ZN(G1347gat));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n651_), .A2(new_n573_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(new_n615_), .A3(new_n644_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n919_), .B1(new_n867_), .B2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n867_), .A2(new_n919_), .A3(new_n922_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(new_n407_), .A3(new_n447_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n867_), .A2(new_n407_), .A3(new_n922_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(G169gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n928_), .A2(new_n932_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n927_), .A2(new_n931_), .A3(new_n933_), .ZN(G1348gat));
  INV_X1    g733(.A(new_n925_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n828_), .B1(new_n935_), .B2(new_n923_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n921_), .B1(new_n871_), .B2(new_n830_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n381_), .A2(new_n424_), .ZN(new_n938_));
  AOI22_X1  g737(.A1(new_n936_), .A2(new_n424_), .B1(new_n937_), .B2(new_n938_), .ZN(G1349gat));
  AOI21_X1  g738(.A(G183gat), .B1(new_n937_), .B2(new_n665_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n343_), .A2(new_n433_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n926_), .B2(new_n941_), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n926_), .A2(new_n901_), .A3(new_n428_), .ZN(new_n943_));
  INV_X1    g742(.A(G190gat), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n713_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n943_), .B1(new_n944_), .B2(new_n945_), .ZN(G1351gat));
  NAND2_X1  g745(.A1(new_n906_), .A2(new_n920_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n406_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n410_), .ZN(G1352gat));
  INV_X1    g748(.A(new_n947_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(new_n828_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g751(.A(new_n343_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(KEYINPUT126), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n950_), .A2(new_n954_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n953_), .A2(KEYINPUT126), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n955_), .A2(new_n956_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n957_), .A2(KEYINPUT127), .A3(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(KEYINPUT127), .ZN(new_n960_));
  OR2_X1    g759(.A1(new_n958_), .A2(KEYINPUT127), .ZN(new_n961_));
  OAI211_X1 g760(.A(new_n960_), .B(new_n961_), .C1(new_n955_), .C2(new_n956_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n959_), .A2(new_n962_), .ZN(G1354gat));
  AND3_X1   g762(.A1(new_n950_), .A2(G218gat), .A3(new_n303_), .ZN(new_n964_));
  AOI21_X1  g763(.A(G218gat), .B1(new_n950_), .B2(new_n901_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n964_), .A2(new_n965_), .ZN(G1355gat));
endmodule


