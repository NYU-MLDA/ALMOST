//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204_));
  INV_X1    g003(.A(G1gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(KEYINPUT81), .A2(G8gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT81), .A2(G8gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n204_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n204_), .B(new_n211_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G29gat), .B(G36gat), .Z(new_n216_));
  XOR2_X1   g015(.A(G43gat), .B(G50gat), .Z(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G29gat), .B(G36gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G43gat), .B(G50gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n215_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT85), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n215_), .A2(new_n225_), .A3(new_n222_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n225_), .B1(new_n215_), .B2(new_n222_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n203_), .B(new_n224_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT15), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n222_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n218_), .A2(KEYINPUT15), .A3(new_n221_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(new_n215_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n215_), .A2(new_n222_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT85), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n236_), .B2(new_n226_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n229_), .B1(new_n237_), .B2(new_n203_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G113gat), .B(G141gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G169gat), .B(G197gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  OR2_X1    g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(KEYINPUT86), .A3(new_n241_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT86), .B1(new_n238_), .B2(new_n241_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n242_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G183gat), .ZN(new_n248_));
  INV_X1    g047(.A(G190gat), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n248_), .A2(new_n249_), .A3(KEYINPUT23), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT23), .B1(new_n248_), .B2(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(G183gat), .B2(G190gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(G169gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n252_), .B(KEYINPUT87), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(new_n250_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G169gat), .B(G176gat), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT24), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT25), .B(G183gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n261_), .B(new_n264_), .C1(KEYINPUT24), .C2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n257_), .B1(new_n259_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G71gat), .B(G99gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(G43gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n267_), .B(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G127gat), .B(G134gat), .Z(new_n271_));
  XOR2_X1   g070(.A(G113gat), .B(G120gat), .Z(new_n272_));
  XOR2_X1   g071(.A(new_n271_), .B(new_n272_), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n270_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275_));
  INV_X1    g074(.A(G15gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT30), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT31), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n279_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n256_), .B1(new_n259_), .B2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(new_n265_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n260_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n286_), .A2(new_n253_), .A3(new_n264_), .A4(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290_));
  INV_X1    g089(.A(G197gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G204gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT92), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G197gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT21), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT91), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n300_), .A2(new_n301_), .ZN(new_n303_));
  OAI221_X1 g102(.A(new_n290_), .B1(KEYINPUT21), .B2(new_n298_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n290_), .A2(new_n299_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n298_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n289_), .A2(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n308_), .B(KEYINPUT20), .C1(new_n307_), .C2(new_n267_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT19), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT96), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n304_), .A2(new_n306_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(new_n284_), .A3(new_n288_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n307_), .A2(new_n267_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n315_), .A2(KEYINPUT20), .A3(new_n316_), .A4(new_n311_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G8gat), .B(G36gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT18), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G64gat), .B(G92gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT32), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n313_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n315_), .A2(KEYINPUT20), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n311_), .B1(new_n324_), .B2(new_n316_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n309_), .A2(new_n312_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT3), .Z(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n333_), .B(KEYINPUT2), .Z(new_n334_));
  OAI211_X1 g133(.A(new_n328_), .B(new_n330_), .C1(new_n332_), .C2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n329_), .B1(KEYINPUT1), .B2(new_n328_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(KEYINPUT1), .B2(new_n328_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n331_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n333_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n340_), .A2(new_n273_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n273_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n341_), .A2(KEYINPUT4), .A3(new_n342_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT100), .ZN(new_n348_));
  INV_X1    g147(.A(new_n342_), .ZN(new_n349_));
  XOR2_X1   g148(.A(KEYINPUT99), .B(KEYINPUT4), .Z(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n342_), .A2(KEYINPUT100), .A3(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n347_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n346_), .B1(new_n354_), .B2(new_n345_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G85gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT0), .B(G57gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n354_), .A2(new_n345_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n346_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n360_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OAI221_X1 g163(.A(new_n323_), .B1(new_n327_), .B2(new_n322_), .C1(new_n361_), .C2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT101), .B1(new_n364_), .B2(KEYINPUT33), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT101), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT33), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n367_), .B(new_n368_), .C1(new_n355_), .C2(new_n360_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n313_), .A2(new_n317_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n321_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT98), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n313_), .A2(new_n317_), .A3(new_n321_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n366_), .A2(new_n369_), .A3(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n354_), .A2(new_n345_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n359_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n364_), .A2(KEYINPUT33), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n374_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n321_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT98), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n365_), .B1(new_n376_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT95), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n335_), .A2(new_n339_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G22gat), .B(G50gat), .Z(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n340_), .A2(KEYINPUT29), .ZN(new_n393_));
  INV_X1    g192(.A(new_n391_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n387_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n391_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n394_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n386_), .A3(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n396_), .A2(KEYINPUT89), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT89), .B1(new_n396_), .B2(new_n399_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n403_), .B(KEYINPUT90), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n405_), .A2(KEYINPUT93), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n388_), .A2(new_n389_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(new_n314_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G78gat), .ZN(new_n409_));
  INV_X1    g208(.A(G78gat), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n410_), .B(new_n406_), .C1(new_n407_), .C2(new_n314_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n405_), .A2(KEYINPUT93), .ZN(new_n412_));
  INV_X1    g211(.A(G106gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n409_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n402_), .B(KEYINPUT94), .C1(new_n415_), .C2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n415_), .A2(new_n416_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n396_), .A2(new_n399_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n418_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT94), .B1(new_n422_), .B2(new_n402_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n385_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n425_));
  INV_X1    g224(.A(new_n402_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n425_), .B1(new_n426_), .B2(new_n418_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n427_), .A2(KEYINPUT95), .A3(new_n420_), .A4(new_n417_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n384_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT27), .B(new_n374_), .C1(new_n327_), .C2(new_n321_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n361_), .A2(new_n364_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n372_), .A2(new_n374_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT102), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT102), .ZN(new_n435_));
  AOI211_X1 g234(.A(new_n435_), .B(KEYINPUT27), .C1(new_n372_), .C2(new_n374_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n430_), .B(new_n431_), .C1(new_n434_), .C2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n282_), .B1(new_n429_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n430_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT103), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT103), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n442_), .B(new_n430_), .C1(new_n434_), .C2(new_n436_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n424_), .A2(new_n428_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n282_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n431_), .A4(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n247_), .B1(new_n439_), .B2(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(G230gat), .A2(G233gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT10), .B(G99gat), .Z(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n413_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G85gat), .B(G92gat), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT9), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT6), .ZN(new_n455_));
  INV_X1    g254(.A(G85gat), .ZN(new_n456_));
  INV_X1    g255(.A(G92gat), .ZN(new_n457_));
  OR3_X1    g256(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT9), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n451_), .A2(new_n453_), .A3(new_n455_), .A4(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G99gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n413_), .A3(KEYINPUT65), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT65), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(G99gat), .B2(G106gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT7), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT66), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT7), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n462_), .A2(new_n464_), .A3(new_n466_), .A4(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT64), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(KEYINPUT64), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n454_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT68), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n477_), .A2(KEYINPUT6), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n479_), .A2(KEYINPUT68), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n476_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(KEYINPUT68), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(KEYINPUT6), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n483_), .A3(new_n454_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n452_), .B1(new_n475_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT69), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n474_), .A2(new_n469_), .A3(new_n481_), .A4(new_n484_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT69), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n452_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n487_), .A2(KEYINPUT8), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n452_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n469_), .A2(new_n474_), .A3(new_n455_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT67), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n474_), .A2(new_n469_), .A3(new_n455_), .A4(KEYINPUT67), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n493_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n460_), .B1(new_n491_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G57gat), .B(G64gat), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n501_), .A2(KEYINPUT11), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(KEYINPUT11), .ZN(new_n503_));
  XOR2_X1   g302(.A(G71gat), .B(G78gat), .Z(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n503_), .A2(new_n504_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n500_), .A2(KEYINPUT70), .A3(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n508_), .B1(new_n507_), .B2(new_n500_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT70), .B1(new_n500_), .B2(new_n507_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n449_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n500_), .B2(new_n507_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n449_), .B1(new_n500_), .B2(new_n507_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n459_), .A2(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n455_), .A2(new_n458_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n517_), .A2(KEYINPUT71), .A3(new_n451_), .A4(new_n453_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n490_), .A2(KEYINPUT8), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n489_), .B1(new_n488_), .B2(new_n452_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n520_), .B1(new_n523_), .B2(new_n498_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n507_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT12), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n513_), .A2(new_n514_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n511_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT72), .ZN(new_n531_));
  XOR2_X1   g330(.A(G176gat), .B(G204gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT74), .ZN(new_n533_));
  XOR2_X1   g332(.A(G120gat), .B(G148gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n530_), .A2(new_n531_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n511_), .B(new_n529_), .C1(KEYINPUT72), .C2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT13), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT13), .B1(new_n538_), .B2(new_n540_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G127gat), .B(G155gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT16), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G183gat), .B(G211gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT84), .B1(new_n549_), .B2(KEYINPUT17), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(new_n215_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(new_n507_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n549_), .A2(KEYINPUT17), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n555_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT77), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT35), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n519_), .B1(new_n491_), .B2(new_n499_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n233_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n222_), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n576_), .B(new_n460_), .C1(new_n491_), .C2(new_n499_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT76), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n571_), .A2(new_n572_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n233_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n524_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n500_), .A2(new_n222_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT76), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .A4(new_n573_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n578_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n579_), .B1(new_n578_), .B2(new_n584_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n567_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n579_), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n524_), .A2(new_n580_), .B1(new_n572_), .B2(new_n571_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n583_), .B1(new_n589_), .B2(new_n582_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n575_), .A2(KEYINPUT76), .A3(new_n577_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n588_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n578_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n564_), .B(KEYINPUT36), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n587_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT80), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT80), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n587_), .A2(new_n595_), .A3(new_n599_), .A4(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n594_), .B(KEYINPUT78), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n592_), .A2(new_n593_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n587_), .A2(new_n603_), .A3(KEYINPUT79), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n604_), .B(KEYINPUT37), .C1(KEYINPUT79), .C2(new_n603_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n560_), .B1(new_n601_), .B2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n448_), .A2(new_n545_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n431_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n205_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n587_), .A2(new_n595_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n439_), .B2(new_n447_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n545_), .A2(new_n246_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT104), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n545_), .A2(KEYINPUT104), .A3(new_n246_), .ZN(new_n618_));
  AND4_X1   g417(.A1(new_n559_), .A2(new_n614_), .A3(new_n617_), .A4(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n608_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(G1gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n609_), .A2(new_n610_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT105), .Z(G1324gat));
  INV_X1    g423(.A(new_n444_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n607_), .A2(new_n625_), .A3(new_n206_), .A4(new_n207_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n619_), .A2(new_n625_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(new_n628_), .A3(G8gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n627_), .B2(G8gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT40), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1325gat));
  NAND3_X1  g432(.A1(new_n607_), .A2(new_n276_), .A3(new_n446_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n619_), .A2(new_n446_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n635_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT41), .B1(new_n635_), .B2(G15gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(G1326gat));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  INV_X1    g438(.A(new_n445_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n607_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n619_), .A2(new_n640_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(G22gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n643_), .A2(new_n644_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n641_), .B1(new_n645_), .B2(new_n646_), .ZN(G1327gat));
  NOR2_X1   g446(.A1(new_n559_), .A2(new_n612_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n545_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n448_), .A2(new_n649_), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n650_), .A2(G29gat), .A3(new_n431_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n617_), .A2(new_n560_), .A3(new_n618_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n439_), .A2(new_n447_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n601_), .A2(new_n605_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n654_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n653_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT44), .B(new_n653_), .C1(new_n658_), .C2(new_n660_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n608_), .A3(new_n664_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n665_), .A2(KEYINPUT108), .A3(G29gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT108), .B1(new_n665_), .B2(G29gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n651_), .B1(new_n666_), .B2(new_n667_), .ZN(G1328gat));
  NOR3_X1   g467(.A1(new_n650_), .A2(G36gat), .A3(new_n444_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n654_), .A2(new_n656_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n659_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n654_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT44), .B1(new_n676_), .B2(new_n653_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n664_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n677_), .A2(new_n678_), .A3(new_n444_), .ZN(new_n679_));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n671_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n671_), .B(new_n682_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1329gat));
  INV_X1    g485(.A(G43gat), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n282_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n663_), .A2(new_n664_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT111), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n663_), .A2(new_n691_), .A3(new_n664_), .A4(new_n688_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n687_), .B1(new_n650_), .B2(new_n282_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n690_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT47), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n690_), .A2(new_n696_), .A3(new_n692_), .A4(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1330gat));
  INV_X1    g497(.A(new_n650_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G50gat), .B1(new_n699_), .B2(new_n640_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n677_), .A2(new_n678_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n640_), .A2(G50gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(G1331gat));
  AOI21_X1  g502(.A(new_n246_), .B1(new_n439_), .B2(new_n447_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n545_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n606_), .ZN(new_n706_));
  INV_X1    g505(.A(G57gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n608_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n614_), .A2(new_n247_), .A3(new_n705_), .A4(new_n559_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G57gat), .B1(new_n709_), .B2(new_n431_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1332gat));
  OAI21_X1  g510(.A(G64gat), .B1(new_n709_), .B2(new_n444_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT48), .ZN(new_n713_));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n706_), .A2(new_n714_), .A3(new_n625_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(G1333gat));
  OAI21_X1  g517(.A(G71gat), .B1(new_n709_), .B2(new_n282_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT49), .ZN(new_n720_));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n706_), .A2(new_n721_), .A3(new_n446_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1334gat));
  OAI21_X1  g522(.A(G78gat), .B1(new_n709_), .B2(new_n445_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT50), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n706_), .A2(new_n410_), .A3(new_n640_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1335gat));
  NAND3_X1  g526(.A1(new_n704_), .A2(new_n705_), .A3(new_n648_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(new_n456_), .A3(new_n608_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n560_), .A2(new_n247_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n676_), .A2(new_n705_), .A3(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(KEYINPUT113), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(KEYINPUT113), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n431_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n730_), .B1(new_n736_), .B2(new_n456_), .ZN(G1336gat));
  NAND3_X1  g536(.A1(new_n729_), .A2(new_n457_), .A3(new_n625_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n734_), .A2(new_n735_), .A3(new_n444_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n457_), .ZN(G1337gat));
  OAI21_X1  g539(.A(G99gat), .B1(new_n733_), .B2(new_n282_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n729_), .A2(new_n446_), .A3(new_n450_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(G1338gat));
  NAND3_X1  g544(.A1(new_n729_), .A2(new_n413_), .A3(new_n640_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n676_), .A2(new_n640_), .A3(new_n705_), .A4(new_n732_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(G106gat), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n747_), .B2(G106gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT53), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n753_), .B(new_n746_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1339gat));
  INV_X1    g554(.A(G113gat), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n237_), .A2(new_n203_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n241_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n223_), .B1(new_n236_), .B2(new_n226_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(new_n203_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n757_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n245_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n243_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n511_), .A2(new_n529_), .A3(new_n539_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n529_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n500_), .A2(new_n507_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n513_), .A2(new_n528_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n449_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT55), .A4(new_n528_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n767_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n537_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT56), .B1(new_n772_), .B2(new_n537_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n765_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT58), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n765_), .B(KEYINPUT58), .C1(new_n773_), .C2(new_n774_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n601_), .A2(new_n777_), .A3(new_n605_), .A4(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n763_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n540_), .B2(new_n538_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782_));
  AOI22_X1  g581(.A1(new_n766_), .A2(new_n529_), .B1(new_n769_), .B2(new_n449_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n539_), .B1(new_n783_), .B2(new_n771_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n784_), .B2(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n774_), .A2(KEYINPUT117), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n537_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n764_), .A2(new_n246_), .A3(KEYINPUT116), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT116), .B1(new_n764_), .B2(new_n246_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n781_), .B1(new_n788_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT57), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n613_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n779_), .B1(new_n792_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n787_), .B1(new_n774_), .B2(KEYINPUT117), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n784_), .A2(new_n782_), .A3(KEYINPUT56), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n791_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n781_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT57), .B1(new_n801_), .B2(new_n612_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT118), .B1(new_n796_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n793_), .B1(new_n792_), .B2(new_n613_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n794_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .A4(new_n779_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n803_), .A2(new_n560_), .A3(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n655_), .A2(new_n247_), .A3(new_n545_), .A4(new_n559_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT54), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n606_), .A2(new_n811_), .A3(new_n247_), .A4(new_n545_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n808_), .A2(new_n813_), .ZN(new_n814_));
  NOR4_X1   g613(.A1(new_n625_), .A2(new_n640_), .A3(new_n431_), .A4(new_n282_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n560_), .B1(new_n796_), .B2(new_n802_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n804_), .A2(new_n805_), .A3(new_n779_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(KEYINPUT119), .A3(new_n560_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n813_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n815_), .A2(new_n823_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n816_), .A2(KEYINPUT59), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n756_), .B1(new_n825_), .B2(new_n246_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n816_), .A2(G113gat), .A3(new_n247_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT120), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n822_), .A2(new_n824_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n246_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G113gat), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  INV_X1    g632(.A(new_n827_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n828_), .A2(new_n835_), .ZN(G1340gat));
  INV_X1    g635(.A(new_n825_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G120gat), .B1(new_n837_), .B2(new_n545_), .ZN(new_n838_));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n545_), .B2(KEYINPUT60), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(KEYINPUT60), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(KEYINPUT121), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(KEYINPUT121), .B2(new_n840_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n838_), .B1(new_n816_), .B2(new_n843_), .ZN(G1341gat));
  NAND2_X1  g643(.A1(new_n559_), .A2(G127gat), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT122), .Z(new_n846_));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n814_), .A2(new_n559_), .A3(new_n815_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n825_), .A2(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(G1342gat));
  OAI21_X1  g648(.A(G134gat), .B1(new_n837_), .B2(new_n655_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n612_), .A2(G134gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n816_), .B2(new_n851_), .ZN(G1343gat));
  AND2_X1   g651(.A1(new_n810_), .A2(new_n812_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n559_), .B1(new_n820_), .B2(KEYINPUT118), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n807_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n445_), .A2(new_n431_), .A3(new_n446_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n444_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT123), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859_));
  INV_X1    g658(.A(new_n857_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n814_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n246_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n705_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g665(.A(KEYINPUT61), .B(G155gat), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n862_), .B2(new_n559_), .ZN(new_n870_));
  AOI211_X1 g669(.A(KEYINPUT124), .B(new_n560_), .C1(new_n858_), .C2(new_n861_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n868_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n859_), .B1(new_n814_), .B2(new_n860_), .ZN(new_n873_));
  AOI211_X1 g672(.A(KEYINPUT123), .B(new_n857_), .C1(new_n808_), .C2(new_n813_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n559_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n862_), .A2(new_n869_), .A3(new_n559_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n867_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n872_), .A2(new_n878_), .ZN(G1346gat));
  NOR2_X1   g678(.A1(new_n873_), .A2(new_n874_), .ZN(new_n880_));
  INV_X1    g679(.A(G162gat), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n880_), .A2(new_n881_), .A3(new_n655_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n612_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(G162gat), .ZN(new_n885_));
  OAI211_X1 g684(.A(KEYINPUT125), .B(new_n881_), .C1(new_n880_), .C2(new_n612_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n882_), .B1(new_n885_), .B2(new_n886_), .ZN(G1347gat));
  AND2_X1   g686(.A1(new_n822_), .A2(new_n445_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n444_), .A2(new_n608_), .A3(new_n282_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n246_), .A3(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT62), .B1(new_n890_), .B2(KEYINPUT22), .ZN(new_n891_));
  OAI21_X1  g690(.A(G169gat), .B1(new_n890_), .B2(KEYINPUT62), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(KEYINPUT62), .B(G169gat), .C1(new_n890_), .C2(KEYINPUT22), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1348gat));
  NAND2_X1  g694(.A1(new_n814_), .A2(new_n445_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n889_), .A2(G176gat), .A3(new_n705_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n888_), .A2(new_n705_), .A3(new_n889_), .ZN(new_n899_));
  INV_X1    g698(.A(G176gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(G1349gat));
  NAND2_X1  g700(.A1(new_n889_), .A2(new_n559_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n896_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n262_), .ZN(new_n904_));
  AOI22_X1  g703(.A1(new_n903_), .A2(new_n248_), .B1(new_n904_), .B2(new_n888_), .ZN(G1350gat));
  NAND4_X1  g704(.A1(new_n888_), .A2(new_n263_), .A3(new_n613_), .A4(new_n889_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n888_), .A2(new_n656_), .A3(new_n889_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n907_), .A2(new_n908_), .A3(G190gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n907_), .B2(G190gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n906_), .B1(new_n909_), .B2(new_n910_), .ZN(G1351gat));
  NOR4_X1   g710(.A1(new_n444_), .A2(new_n445_), .A3(new_n608_), .A4(new_n446_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n814_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n247_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n291_), .ZN(G1352gat));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n545_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n295_), .ZN(G1353gat));
  INV_X1    g716(.A(new_n913_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n559_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  AOI21_X1  g722(.A(G218gat), .B1(new_n918_), .B2(new_n613_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n656_), .A2(G218gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT127), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n918_), .B2(new_n926_), .ZN(G1355gat));
endmodule


