//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n851_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G85gat), .B(G92gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G85gat), .A3(G92gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT8), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT64), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n214_), .A2(new_n216_), .A3(new_n207_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n207_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT65), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n207_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n213_), .A2(KEYINPUT64), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n214_), .A2(new_n216_), .A3(new_n207_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT7), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n219_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n212_), .B1(new_n229_), .B2(new_n205_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n205_), .A2(new_n212_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(new_n228_), .B2(new_n208_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n211_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT66), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G43gat), .B(G50gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G29gat), .B(G36gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT72), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT73), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n236_), .A2(KEYINPUT72), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT73), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(KEYINPUT72), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n235_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n238_), .A2(new_n242_), .A3(new_n235_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n247_), .B(new_n211_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n234_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT15), .ZN(new_n250_));
  INV_X1    g049(.A(new_n245_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(new_n243_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n244_), .A2(KEYINPUT15), .A3(new_n245_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(new_n233_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(KEYINPUT74), .A3(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n249_), .A2(new_n254_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT35), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n249_), .A2(KEYINPUT74), .A3(new_n254_), .A4(new_n258_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n260_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G190gat), .B(G218gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G134gat), .B(G162gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(KEYINPUT36), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n268_), .B(KEYINPUT36), .Z(new_n271_));
  NAND4_X1  g070(.A1(new_n260_), .A2(new_n263_), .A3(new_n264_), .A4(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT75), .B(KEYINPUT37), .Z(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT76), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT37), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT76), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n270_), .A2(new_n278_), .A3(new_n272_), .A4(new_n273_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G71gat), .B(G78gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(G57gat), .B(G64gat), .Z(new_n282_));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G57gat), .B(G64gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT11), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n281_), .A3(KEYINPUT11), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n288_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT77), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G15gat), .B(G22gat), .ZN(new_n298_));
  INV_X1    g097(.A(G1gat), .ZN(new_n299_));
  INV_X1    g098(.A(G8gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT14), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n297_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n297_), .A2(new_n303_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n294_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G127gat), .B(G155gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT16), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G183gat), .B(G211gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT17), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n310_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n297_), .B(new_n302_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n309_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n293_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n315_), .A2(new_n316_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n311_), .A2(new_n318_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n319_), .A2(new_n321_), .A3(KEYINPUT78), .ZN(new_n327_));
  INV_X1    g126(.A(new_n292_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(KEYINPUT69), .A3(new_n290_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n326_), .A2(new_n327_), .A3(new_n329_), .A4(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n317_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n326_), .A2(new_n327_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n324_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT79), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n337_), .B(new_n324_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n280_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n341_), .B(KEYINPUT80), .Z(new_n342_));
  INV_X1    g141(.A(KEYINPUT71), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n234_), .A2(new_n293_), .A3(new_n248_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n233_), .A2(new_n331_), .A3(new_n329_), .A4(KEYINPUT12), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n234_), .A2(new_n248_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n294_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT12), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G230gat), .A2(G233gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n344_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n293_), .B1(new_n234_), .B2(new_n248_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G120gat), .B(G148gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(G176gat), .B(G204gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n353_), .A2(new_n357_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT13), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n363_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n353_), .A2(new_n357_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n362_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT13), .B1(new_n370_), .B2(new_n364_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n343_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n366_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(KEYINPUT13), .A3(new_n364_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(KEYINPUT71), .A3(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G113gat), .B(G141gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G169gat), .B(G197gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n252_), .A2(new_n253_), .A3(new_n306_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n306_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G229gat), .A2(G233gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n385_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n246_), .A2(new_n320_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n383_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT82), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n390_), .A2(KEYINPUT81), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n390_), .B2(KEYINPUT81), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n381_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n390_), .A2(KEYINPUT81), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT82), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n390_), .A2(KEYINPUT81), .A3(new_n391_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n380_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n394_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n377_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G127gat), .B(G134gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT89), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n402_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT88), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G141gat), .A2(G148gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT3), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G141gat), .A2(G148gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT2), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(KEYINPUT1), .B2(new_n413_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(KEYINPUT1), .B2(new_n413_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n408_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n410_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n407_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n405_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n417_), .B(new_n421_), .C1(new_n424_), .C2(new_n403_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT4), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n423_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n426_), .A2(new_n428_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G1gat), .B(G29gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G85gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT0), .B(G57gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n436_), .B(new_n437_), .Z(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n432_), .A2(new_n440_), .A3(new_n433_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n441_), .A3(KEYINPUT100), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT100), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n434_), .A2(new_n443_), .A3(new_n438_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G211gat), .B(G218gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT21), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G197gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G204gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n448_), .A2(G204gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n447_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT92), .ZN(new_n456_));
  OR3_X1    g255(.A1(new_n454_), .A2(KEYINPUT91), .A3(KEYINPUT21), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT91), .B1(new_n454_), .B2(KEYINPUT21), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n453_), .A2(new_n449_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT21), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n457_), .A2(new_n458_), .A3(new_n445_), .A4(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G183gat), .ZN(new_n463_));
  INV_X1    g262(.A(G190gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT23), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT23), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(G183gat), .A3(G190gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(G183gat), .B2(G190gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT85), .B(G176gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT22), .B(G169gat), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n470_), .A2(new_n471_), .B1(G169gat), .B2(G176gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(KEYINPUT86), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(new_n465_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G169gat), .A2(G176gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(KEYINPUT24), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n476_), .B(KEYINPUT83), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G169gat), .A2(G176gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(KEYINPUT24), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT25), .B(G183gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT26), .B(G190gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n473_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n462_), .A2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n468_), .B1(new_n479_), .B2(KEYINPUT24), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT84), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n485_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n489_), .B2(new_n485_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n475_), .B1(G183gat), .B2(G190gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n472_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT20), .B(new_n487_), .C1(new_n494_), .C2(new_n462_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G226gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT19), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n462_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n497_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n462_), .A2(new_n486_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n499_), .A2(KEYINPUT20), .A3(new_n500_), .A4(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G8gat), .B(G36gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT18), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G64gat), .B(G92gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT32), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n498_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n442_), .A2(new_n444_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n501_), .A2(KEYINPUT99), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n499_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT99), .B1(new_n501_), .B2(new_n510_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n497_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n495_), .A2(new_n497_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n507_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n498_), .A2(new_n506_), .A3(new_n502_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT97), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT97), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n498_), .A2(new_n502_), .A3(new_n519_), .A4(new_n506_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n498_), .A2(new_n502_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n506_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n518_), .A2(new_n520_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n440_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT33), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT33), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n427_), .A2(new_n431_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n428_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n426_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n438_), .B1(new_n530_), .B2(new_n429_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n526_), .B1(new_n532_), .B2(new_n525_), .ZN(new_n533_));
  OAI22_X1  g332(.A1(new_n509_), .A2(new_n516_), .B1(new_n524_), .B2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n422_), .A2(KEYINPUT29), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT28), .Z(new_n536_));
  XNOR2_X1  g335(.A(G22gat), .B(G50gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n422_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT94), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n422_), .A2(new_n542_), .A3(new_n539_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n462_), .A3(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(G228gat), .A3(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G78gat), .B(G106gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n422_), .A2(KEYINPUT29), .B1(G228gat), .B2(G233gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n462_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n538_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n547_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n550_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n545_), .A2(KEYINPUT95), .A3(new_n547_), .A4(new_n549_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n538_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n554_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AOI211_X1 g359(.A(KEYINPUT96), .B(new_n538_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n534_), .B(new_n553_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n553_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n442_), .A2(new_n444_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n514_), .A2(new_n515_), .ZN(new_n566_));
  OAI211_X1 g365(.A(KEYINPUT27), .B(new_n517_), .C1(new_n566_), .C2(new_n506_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT27), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n524_), .A2(KEYINPUT101), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT101), .B1(new_n524_), .B2(new_n568_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n567_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n562_), .B1(new_n565_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G227gat), .A2(G233gat), .ZN(new_n573_));
  INV_X1    g372(.A(G15gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT30), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n494_), .B(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n407_), .B(KEYINPUT31), .Z(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT87), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n577_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G71gat), .B(G99gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(G43gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n580_), .B(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n571_), .A2(new_n563_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n564_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n572_), .A2(new_n583_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n342_), .A2(new_n400_), .A3(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n299_), .A3(new_n585_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT38), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT103), .Z(new_n593_));
  INV_X1    g392(.A(new_n276_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n587_), .A2(new_n594_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n377_), .A2(new_n335_), .A3(new_n399_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n299_), .B1(new_n597_), .B2(new_n585_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT102), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n593_), .B(new_n599_), .C1(new_n591_), .C2(new_n590_), .ZN(G1324gat));
  NAND3_X1  g399(.A1(new_n589_), .A2(new_n300_), .A3(new_n571_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT104), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n597_), .A2(new_n571_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n606_), .B2(G8gat), .ZN(new_n607_));
  AOI211_X1 g406(.A(KEYINPUT39), .B(new_n300_), .C1(new_n597_), .C2(new_n571_), .ZN(new_n608_));
  OAI22_X1  g407(.A1(new_n603_), .A2(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT40), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI221_X1 g410(.A(KEYINPUT40), .B1(new_n607_), .B2(new_n608_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1325gat));
  INV_X1    g412(.A(new_n583_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n574_), .B1(new_n597_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n589_), .A2(new_n574_), .A3(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n597_), .B2(new_n563_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n589_), .A2(new_n619_), .A3(new_n563_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1327gat));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n625_), .B1(new_n587_), .B2(new_n280_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n280_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n524_), .A2(new_n568_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n524_), .A2(KEYINPUT101), .A3(new_n568_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n632_), .A2(new_n567_), .A3(new_n564_), .A4(new_n563_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n614_), .B1(new_n633_), .B2(new_n562_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n586_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n635_), .A2(new_n571_), .A3(new_n563_), .ZN(new_n636_));
  OAI211_X1 g435(.A(KEYINPUT43), .B(new_n627_), .C1(new_n634_), .C2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n626_), .A2(new_n339_), .A3(new_n400_), .A4(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n627_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n340_), .B1(new_n641_), .B2(new_n625_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n642_), .A2(KEYINPUT44), .A3(new_n400_), .A4(new_n637_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n640_), .A2(new_n643_), .A3(G29gat), .A4(new_n585_), .ZN(new_n644_));
  INV_X1    g443(.A(G29gat), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n340_), .A2(new_n276_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n588_), .A2(new_n400_), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(new_n647_), .B2(new_n564_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n644_), .A2(new_n648_), .ZN(G1328gat));
  NAND3_X1  g448(.A1(new_n640_), .A2(new_n571_), .A3(new_n643_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G36gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n571_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(G36gat), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n588_), .A2(new_n400_), .A3(new_n646_), .A4(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT45), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n651_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT46), .B1(new_n658_), .B2(KEYINPUT106), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n660_), .B(new_n661_), .C1(new_n651_), .C2(new_n657_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n659_), .A2(new_n662_), .ZN(G1329gat));
  NAND4_X1  g462(.A1(new_n640_), .A2(new_n643_), .A3(G43gat), .A4(new_n614_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n647_), .A2(new_n583_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(G43gat), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g466(.A1(new_n640_), .A2(new_n643_), .A3(G50gat), .A4(new_n563_), .ZN(new_n668_));
  INV_X1    g467(.A(G50gat), .ZN(new_n669_));
  INV_X1    g468(.A(new_n563_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n647_), .B2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n668_), .A2(new_n671_), .ZN(G1331gat));
  AOI21_X1  g471(.A(new_n339_), .B1(new_n398_), .B2(new_n394_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n595_), .A2(new_n377_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n675_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(G57gat), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n564_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n399_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n587_), .A2(new_n682_), .A3(new_n376_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n342_), .A3(new_n585_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(KEYINPUT107), .A3(new_n679_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT107), .B1(new_n684_), .B2(new_n679_), .ZN(new_n687_));
  OAI22_X1  g486(.A1(new_n678_), .A2(new_n681_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n688_), .A2(KEYINPUT109), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(KEYINPUT109), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1332gat));
  NAND2_X1  g490(.A1(new_n683_), .A2(new_n342_), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n692_), .A2(G64gat), .A3(new_n652_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n676_), .A2(new_n571_), .A3(new_n677_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(new_n695_), .A3(G64gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n694_), .B2(G64gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(G1333gat));
  NAND3_X1  g497(.A1(new_n676_), .A2(new_n614_), .A3(new_n677_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT49), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(G71gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(G71gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n583_), .A2(G71gat), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT110), .Z(new_n704_));
  OAI22_X1  g503(.A1(new_n701_), .A2(new_n702_), .B1(new_n692_), .B2(new_n704_), .ZN(G1334gat));
  OR3_X1    g504(.A1(new_n692_), .A2(G78gat), .A3(new_n670_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n676_), .A2(new_n563_), .A3(new_n677_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT50), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(G78gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n707_), .B2(G78gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n587_), .A2(new_n682_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(new_n377_), .A3(new_n646_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n585_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT111), .Z(new_n716_));
  NOR2_X1   g515(.A1(new_n376_), .A2(new_n682_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n626_), .A2(new_n339_), .A3(new_n637_), .A4(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n719_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n720_), .A2(G85gat), .A3(new_n585_), .A4(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n716_), .A2(new_n722_), .ZN(G1336gat));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n571_), .A3(new_n721_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G92gat), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n652_), .A2(G92gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n713_), .B2(new_n726_), .ZN(G1337gat));
  NAND3_X1  g526(.A1(new_n714_), .A2(new_n202_), .A3(new_n614_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G99gat), .B1(new_n718_), .B2(new_n583_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n728_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n731_), .B(new_n732_), .Z(G1338gat));
  NOR3_X1   g532(.A1(new_n713_), .A2(G106gat), .A3(new_n670_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n203_), .B1(new_n735_), .B2(KEYINPUT52), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n718_), .B2(new_n670_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n735_), .B2(KEYINPUT52), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n735_), .A2(KEYINPUT52), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n736_), .B(new_n739_), .C1(new_n718_), .C2(new_n670_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n734_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n741_), .B(new_n743_), .ZN(G1339gat));
  INV_X1    g543(.A(new_n335_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n394_), .A2(new_n398_), .A3(new_n364_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT12), .B1(new_n348_), .B2(new_n294_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n354_), .B1(new_n747_), .B2(new_n346_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT117), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n344_), .B(new_n345_), .C1(new_n356_), .C2(KEYINPUT12), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n354_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n347_), .A2(new_n351_), .A3(KEYINPUT55), .A4(new_n352_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n754_), .A3(new_n354_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n749_), .A2(new_n752_), .A3(new_n753_), .A4(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n362_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n362_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n746_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n382_), .A2(new_n384_), .A3(new_n387_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n385_), .B1(new_n388_), .B2(new_n383_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n380_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n381_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n370_), .B2(new_n364_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n276_), .B1(new_n761_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT57), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n394_), .A2(new_n398_), .A3(new_n364_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n362_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT56), .B1(new_n756_), .B2(new_n362_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n767_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n276_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n769_), .A2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n365_), .A2(new_n766_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n280_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n759_), .A2(new_n760_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n783_), .A2(KEYINPUT118), .A3(KEYINPUT58), .A4(new_n779_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT58), .B(new_n779_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n782_), .A2(new_n784_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n745_), .B1(new_n778_), .B2(new_n788_), .ZN(new_n789_));
  XOR2_X1   g588(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n790_));
  AND3_X1   g589(.A1(new_n673_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n280_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n791_), .A2(new_n280_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT119), .B1(new_n789_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n776_), .B1(new_n775_), .B2(new_n276_), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT57), .B(new_n594_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n788_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n335_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n795_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NOR4_X1   g602(.A1(new_n571_), .A2(new_n564_), .A3(new_n563_), .A4(new_n583_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n796_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(G113gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n682_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n795_), .B1(new_n799_), .B2(new_n339_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n804_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT120), .B1(new_n809_), .B2(new_n813_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n805_), .A2(KEYINPUT59), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n817_), .A2(new_n682_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n808_), .B1(new_n818_), .B2(new_n807_), .ZN(G1340gat));
  INV_X1    g618(.A(G120gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n376_), .B2(KEYINPUT60), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(KEYINPUT60), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(KEYINPUT121), .B2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n806_), .B(new_n823_), .C1(KEYINPUT121), .C2(new_n821_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n817_), .A2(new_n377_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n820_), .ZN(G1341gat));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n806_), .A2(new_n827_), .A3(new_n340_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n817_), .A2(new_n745_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n827_), .ZN(G1342gat));
  AOI21_X1  g629(.A(G134gat), .B1(new_n806_), .B2(new_n594_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT122), .B(G134gat), .Z(new_n832_));
  NOR2_X1   g631(.A1(new_n280_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n831_), .B1(new_n817_), .B2(new_n833_), .ZN(G1343gat));
  AOI21_X1  g633(.A(new_n802_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n835_));
  AOI211_X1 g634(.A(KEYINPUT119), .B(new_n795_), .C1(new_n799_), .C2(new_n335_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n670_), .A2(new_n614_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n839_), .A2(new_n571_), .A3(new_n564_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT123), .B1(new_n837_), .B2(new_n840_), .ZN(new_n841_));
  AND4_X1   g640(.A1(KEYINPUT123), .A2(new_n796_), .A3(new_n803_), .A4(new_n840_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n682_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G141gat), .ZN(new_n844_));
  INV_X1    g643(.A(G141gat), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n845_), .B(new_n682_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1344gat));
  OAI21_X1  g646(.A(new_n377_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G148gat), .ZN(new_n849_));
  INV_X1    g648(.A(G148gat), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n850_), .B(new_n377_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1345gat));
  OAI21_X1  g651(.A(new_n340_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n854_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n340_), .B(new_n856_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1346gat));
  INV_X1    g657(.A(G162gat), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n859_), .B(new_n594_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n837_), .A2(KEYINPUT123), .A3(new_n840_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n796_), .A2(new_n803_), .A3(new_n840_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n280_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n860_), .B1(new_n859_), .B2(new_n865_), .ZN(G1347gat));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n652_), .A2(new_n563_), .A3(new_n635_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n810_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n399_), .ZN(new_n871_));
  INV_X1    g670(.A(G169gat), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n867_), .B(new_n868_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n874_));
  OAI221_X1 g673(.A(new_n874_), .B1(KEYINPUT124), .B2(KEYINPUT62), .C1(new_n870_), .C2(new_n399_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n471_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n875_), .A3(new_n876_), .ZN(G1348gat));
  INV_X1    g676(.A(new_n870_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n377_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n835_), .A2(new_n836_), .A3(new_n563_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n652_), .A2(new_n635_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n377_), .A2(new_n881_), .A3(G176gat), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n879_), .A2(new_n470_), .B1(new_n880_), .B2(new_n882_), .ZN(G1349gat));
  NOR3_X1   g682(.A1(new_n870_), .A2(new_n335_), .A3(new_n482_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(new_n340_), .A3(new_n881_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n463_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n870_), .B2(new_n280_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n594_), .A2(new_n483_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n870_), .B2(new_n888_), .ZN(G1351gat));
  NOR3_X1   g688(.A1(new_n839_), .A2(new_n652_), .A3(new_n585_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n837_), .A2(new_n682_), .A3(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g691(.A1(new_n837_), .A2(new_n377_), .A3(new_n890_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n837_), .A2(new_n745_), .A3(new_n890_), .A4(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  XOR2_X1   g696(.A(new_n897_), .B(KEYINPUT125), .Z(new_n898_));
  XNOR2_X1  g697(.A(new_n896_), .B(new_n898_), .ZN(G1354gat));
  AND2_X1   g698(.A1(new_n837_), .A2(new_n890_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n594_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT126), .B(G218gat), .Z(new_n902_));
  NOR2_X1   g701(.A1(new_n280_), .A2(new_n902_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n901_), .A2(new_n902_), .B1(new_n900_), .B2(new_n903_), .ZN(G1355gat));
endmodule


