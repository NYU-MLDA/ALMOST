//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G43gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G227gat), .A2(G233gat), .ZN(new_n204_));
  INV_X1    g003(.A(G15gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n203_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(G190gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT23), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT81), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT79), .B(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n218_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OR3_X1    g022(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT80), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n217_), .A2(new_n223_), .A3(new_n224_), .A4(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT22), .ZN(new_n231_));
  OAI21_X1  g030(.A(G169gat), .B1(new_n231_), .B2(KEYINPUT83), .ZN(new_n232_));
  INV_X1    g031(.A(G176gat), .ZN(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT22), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n232_), .B(new_n233_), .C1(KEYINPUT83), .C2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n219_), .A2(new_n209_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT84), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n211_), .A2(new_n214_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n226_), .B(new_n236_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n230_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT30), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n208_), .B1(new_n245_), .B2(KEYINPUT85), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT85), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n246_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G127gat), .B(G134gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G113gat), .B(G120gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n250_), .B(new_n251_), .Z(new_n252_));
  OR2_X1    g051(.A1(new_n252_), .A2(KEYINPUT31), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(KEYINPUT31), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n253_), .A2(KEYINPUT86), .A3(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n249_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G8gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G64gat), .B(G92gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G197gat), .B(G204gat), .Z(new_n262_));
  INV_X1    g061(.A(KEYINPUT93), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT21), .ZN(new_n264_));
  XOR2_X1   g063(.A(G211gat), .B(G218gat), .Z(new_n265_));
  OR2_X1    g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n265_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n262_), .A2(KEYINPUT21), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n230_), .A3(new_n242_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n231_), .A2(G169gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n235_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n226_), .B1(G176gat), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n209_), .A2(new_n210_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n217_), .B2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n227_), .B1(G169gat), .B2(G176gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n239_), .A2(new_n224_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G190gat), .ZN(new_n278_));
  AOI211_X1 g077(.A(new_n276_), .B(new_n277_), .C1(new_n218_), .C2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n270_), .B(KEYINPUT20), .C1(new_n280_), .C2(new_n269_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT98), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT19), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n269_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n269_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n243_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n284_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n286_), .A2(new_n288_), .A3(KEYINPUT20), .A4(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n282_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n261_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n281_), .A2(new_n284_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT98), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n295_), .A2(new_n260_), .A3(new_n290_), .A4(new_n285_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(KEYINPUT99), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n295_), .A2(new_n290_), .A3(new_n285_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT99), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n261_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n297_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n286_), .A2(KEYINPUT20), .A3(new_n288_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n284_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n284_), .B2(new_n281_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n261_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(KEYINPUT27), .A3(new_n296_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G78gat), .B(G106gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT95), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(KEYINPUT97), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT90), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n313_), .B(new_n316_), .C1(KEYINPUT3), .C2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(KEYINPUT87), .Z(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n319_), .B(KEYINPUT88), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n321_), .A2(KEYINPUT1), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n323_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n330_));
  XOR2_X1   g129(.A(G141gat), .B(G148gat), .Z(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n330_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n324_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n269_), .B1(new_n335_), .B2(KEYINPUT29), .ZN(new_n336_));
  AND2_X1   g135(.A1(KEYINPUT92), .A2(G228gat), .ZN(new_n337_));
  NOR2_X1   g136(.A1(KEYINPUT92), .A2(G228gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(G233gat), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT94), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n336_), .A2(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(KEYINPUT94), .B(G233gat), .C1(new_n337_), .C2(new_n338_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n318_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n329_), .A2(new_n331_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT89), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n345_), .B2(new_n332_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n287_), .B(new_n342_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n311_), .B1(new_n341_), .B2(new_n349_), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n341_), .A2(new_n349_), .A3(new_n311_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT28), .B1(new_n335_), .B2(KEYINPUT29), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT91), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT28), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n346_), .A2(new_n354_), .A3(new_n347_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n353_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G22gat), .B(G50gat), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n355_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n354_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT91), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n359_), .B1(new_n364_), .B2(new_n356_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n350_), .B(new_n351_), .C1(new_n361_), .C2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT96), .B1(new_n341_), .B2(new_n349_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT96), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n348_), .B(new_n368_), .C1(new_n336_), .C2(new_n340_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n310_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n364_), .A2(new_n359_), .A3(new_n356_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n369_), .A2(new_n310_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n360_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n366_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n335_), .A2(new_n252_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n252_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n346_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n378_), .A3(KEYINPUT4), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n346_), .A2(KEYINPUT4), .A3(new_n377_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n376_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT100), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n376_), .A2(new_n378_), .A3(KEYINPUT100), .A4(new_n381_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n383_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT0), .B(G57gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n383_), .A2(new_n386_), .A3(new_n392_), .A4(new_n387_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR4_X1   g195(.A1(new_n256_), .A2(new_n308_), .A3(new_n375_), .A4(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n302_), .A2(new_n307_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n396_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n375_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n297_), .A2(new_n301_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n379_), .A2(new_n381_), .A3(new_n380_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n376_), .A2(new_n378_), .A3(new_n382_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n393_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT101), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT101), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n393_), .A4(new_n403_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n395_), .A2(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n386_), .A2(new_n387_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n412_), .A2(KEYINPUT33), .A3(new_n392_), .A4(new_n383_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n401_), .A2(new_n409_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n260_), .A2(KEYINPUT32), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n299_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n416_), .B2(new_n305_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n396_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n414_), .A2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n400_), .B1(new_n420_), .B2(new_n375_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n397_), .B1(new_n421_), .B2(new_n256_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G29gat), .B(G36gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G43gat), .B(G50gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT77), .Z(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT72), .B(G15gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G22gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT73), .B(G1gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT74), .B(G8gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G1gat), .B(G8gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  OR3_X1    g233(.A1(new_n428_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n434_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n426_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n425_), .B(KEYINPUT77), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G229gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n425_), .B(KEYINPUT15), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n438_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G113gat), .B(G141gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G169gat), .B(G197gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n444_), .A2(new_n447_), .A3(new_n451_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n444_), .A2(KEYINPUT78), .A3(new_n447_), .A4(new_n451_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n453_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT66), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G85gat), .A2(G92gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n463_), .A2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n471_));
  NOR2_X1   g270(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n472_));
  OAI22_X1  g271(.A1(new_n471_), .A2(new_n472_), .B1(G99gat), .B2(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT6), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(G99gat), .A3(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n479_));
  INV_X1    g278(.A(G99gat), .ZN(new_n480_));
  INV_X1    g279(.A(G106gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(new_n478_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n470_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT64), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n476_), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n474_), .A2(KEYINPUT6), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n475_), .A2(new_n477_), .A3(KEYINPUT64), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n488_), .A2(new_n473_), .A3(new_n482_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n463_), .A2(new_n469_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(KEYINPUT8), .A2(new_n484_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n475_), .A2(new_n477_), .A3(KEYINPUT64), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT64), .B1(new_n475_), .B2(new_n477_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT10), .B(G99gat), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(G106gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n468_), .A2(KEYINPUT9), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n461_), .A2(new_n462_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(KEYINPUT9), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT67), .B1(new_n494_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n508_));
  XOR2_X1   g307(.A(G71gat), .B(G78gat), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n508_), .A2(new_n509_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT67), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n473_), .A2(new_n482_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n492_), .B1(new_n497_), .B2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n491_), .B1(new_n470_), .B2(new_n483_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n513_), .B(new_n503_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n505_), .A2(new_n512_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n484_), .A2(KEYINPUT8), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n490_), .A2(new_n493_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n503_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n512_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(KEYINPUT12), .A3(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n518_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n513_), .B1(new_n521_), .B2(new_n503_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n517_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n523_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n525_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n528_), .A2(new_n518_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n532_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G120gat), .B(G148gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(KEYINPUT69), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n532_), .B(new_n539_), .C1(new_n533_), .C2(new_n531_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n542_), .A2(KEYINPUT13), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT13), .B1(new_n542_), .B2(new_n543_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n505_), .A2(new_n425_), .A3(new_n517_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n522_), .A2(new_n445_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(KEYINPUT71), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT35), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n554_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n548_), .A2(new_n549_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n557_), .A2(new_n558_), .B1(KEYINPUT36), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n555_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n555_), .A2(new_n566_), .A3(new_n556_), .A4(new_n562_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT37), .ZN(new_n569_));
  XOR2_X1   g368(.A(G127gat), .B(G155gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT76), .ZN(new_n571_));
  XOR2_X1   g370(.A(G183gat), .B(G211gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n575_), .B(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n512_), .B(new_n580_), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(new_n437_), .ZN(new_n582_));
  MUX2_X1   g381(.A(new_n578_), .B(new_n579_), .S(new_n582_), .Z(new_n583_));
  NAND2_X1  g382(.A1(new_n569_), .A2(new_n583_), .ZN(new_n584_));
  NOR4_X1   g383(.A1(new_n422_), .A2(new_n460_), .A3(new_n547_), .A4(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n396_), .A2(KEYINPUT102), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n396_), .A2(KEYINPUT102), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n430_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(KEYINPUT38), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(KEYINPUT38), .ZN(new_n593_));
  INV_X1    g392(.A(new_n568_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n422_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n546_), .A2(new_n459_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n583_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G1gat), .B1(new_n600_), .B2(new_n399_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n592_), .A2(new_n593_), .A3(new_n601_), .ZN(G1324gat));
  XNOR2_X1  g401(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n308_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(G8gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT39), .ZN(new_n606_));
  INV_X1    g405(.A(new_n431_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n585_), .A2(new_n308_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n603_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n605_), .A2(KEYINPUT39), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n604_), .B2(G8gat), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n608_), .B(new_n603_), .C1(new_n610_), .C2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n609_), .A2(new_n614_), .ZN(G1325gat));
  INV_X1    g414(.A(new_n256_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n205_), .B1(new_n599_), .B2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT41), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n585_), .A2(new_n205_), .A3(new_n616_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1326gat));
  INV_X1    g419(.A(G22gat), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n585_), .A2(new_n621_), .A3(new_n375_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n375_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G22gat), .B1(new_n600_), .B2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n624_), .A2(KEYINPUT42), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(KEYINPUT42), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n622_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(KEYINPUT104), .B(new_n622_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1327gat));
  NOR2_X1   g430(.A1(new_n422_), .A2(new_n460_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n568_), .A2(new_n583_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n546_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n396_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT37), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n568_), .B(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n640_), .B2(KEYINPUT105), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n641_), .B1(new_n422_), .B2(new_n569_), .ZN(new_n642_));
  AND4_X1   g441(.A1(new_n375_), .A2(new_n399_), .A3(new_n302_), .A4(new_n307_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n375_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n256_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n256_), .A2(new_n308_), .A3(new_n375_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n399_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n641_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n640_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n642_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n596_), .A2(new_n583_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(KEYINPUT44), .A3(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n588_), .A2(G29gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n637_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  NOR3_X1   g459(.A1(new_n635_), .A2(G36gat), .A3(new_n398_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT45), .Z(new_n662_));
  OAI21_X1  g461(.A(G36gat), .B1(new_n657_), .B2(new_n398_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n662_), .A2(new_n663_), .A3(KEYINPUT46), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  NAND2_X1  g467(.A1(new_n616_), .A2(G43gat), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n635_), .A2(new_n256_), .ZN(new_n670_));
  OAI22_X1  g469(.A1(new_n657_), .A2(new_n669_), .B1(G43gat), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g471(.A(G50gat), .B1(new_n657_), .B2(new_n623_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n623_), .A2(G50gat), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT106), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n635_), .B2(new_n675_), .ZN(G1331gat));
  NOR3_X1   g475(.A1(new_n546_), .A2(new_n459_), .A3(new_n597_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n595_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G57gat), .B1(new_n679_), .B2(new_n399_), .ZN(new_n680_));
  NOR4_X1   g479(.A1(new_n422_), .A2(new_n459_), .A3(new_n546_), .A4(new_n584_), .ZN(new_n681_));
  INV_X1    g480(.A(G57gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n588_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1332gat));
  NOR2_X1   g483(.A1(new_n398_), .A2(G64gat), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT107), .Z(new_n686_));
  NAND2_X1  g485(.A1(new_n681_), .A2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G64gat), .B1(new_n679_), .B2(new_n398_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT48), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT48), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OAI211_X1 g492(.A(KEYINPUT108), .B(new_n687_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1333gat));
  INV_X1    g494(.A(G71gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n678_), .B2(new_n616_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT49), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n681_), .A2(new_n696_), .A3(new_n616_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1334gat));
  INV_X1    g499(.A(G78gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n678_), .B2(new_n375_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT50), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n681_), .A2(new_n701_), .A3(new_n375_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1335gat));
  NOR2_X1   g504(.A1(new_n546_), .A2(new_n459_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n597_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n649_), .B1(new_n648_), .B2(new_n640_), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n569_), .B(new_n641_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n708_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G85gat), .B1(new_n713_), .B2(new_n399_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n648_), .A2(new_n706_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n633_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(new_n464_), .A3(new_n588_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n718_), .ZN(G1336gat));
  NOR3_X1   g518(.A1(new_n713_), .A2(new_n465_), .A3(new_n398_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n465_), .B1(new_n716_), .B2(new_n398_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT110), .Z(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1337gat));
  OR2_X1    g522(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n724_));
  NAND2_X1  g523(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n711_), .B(KEYINPUT109), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n480_), .B1(new_n726_), .B2(new_n616_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n716_), .A2(new_n256_), .A3(new_n498_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n724_), .B(new_n725_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G99gat), .B1(new_n713_), .B2(new_n256_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n728_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n730_), .A2(KEYINPUT111), .A3(KEYINPUT51), .A4(new_n731_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n729_), .A2(new_n732_), .ZN(G1338gat));
  NAND3_X1  g532(.A1(new_n717_), .A2(new_n481_), .A3(new_n375_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n375_), .B(new_n708_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT112), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n651_), .A2(new_n737_), .A3(new_n375_), .A4(new_n708_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  OAI21_X1  g539(.A(G106gat), .B1(new_n740_), .B2(KEYINPUT113), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n739_), .A2(new_n742_), .B1(KEYINPUT113), .B2(new_n740_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(KEYINPUT113), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n744_), .B(new_n741_), .C1(new_n736_), .C2(new_n738_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n734_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n734_), .C1(new_n743_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  NAND2_X1  g549(.A1(new_n646_), .A2(new_n588_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT58), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n512_), .B1(new_n505_), .B2(new_n517_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n518_), .B(new_n524_), .C1(new_n753_), .C2(KEYINPUT12), .ZN(new_n754_));
  INV_X1    g553(.A(new_n531_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT114), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT55), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n532_), .A2(KEYINPUT114), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n531_), .B1(new_n525_), .B2(new_n530_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n757_), .A2(new_n759_), .A3(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT56), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n541_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n454_), .A2(new_n455_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n438_), .A2(new_n443_), .A3(new_n446_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n451_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n765_), .A2(new_n457_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(new_n543_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n764_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n760_), .B1(new_n756_), .B2(KEYINPUT55), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n540_), .B1(new_n771_), .B2(new_n759_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n763_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n752_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n762_), .A2(new_n541_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT56), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n776_), .A2(KEYINPUT58), .A3(new_n764_), .A4(new_n769_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n640_), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n763_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n459_), .A2(new_n543_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n542_), .A2(new_n543_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n768_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n594_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n778_), .B1(new_n786_), .B2(KEYINPUT57), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n788_), .B(new_n594_), .C1(new_n783_), .C2(new_n785_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n597_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n569_), .A2(new_n546_), .A3(new_n460_), .A4(new_n583_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n751_), .B1(new_n790_), .B2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(G113gat), .B1(new_n795_), .B2(new_n459_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT116), .Z(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  INV_X1    g597(.A(new_n751_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n780_), .B1(new_n762_), .B2(new_n541_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n782_), .B1(new_n800_), .B2(KEYINPUT56), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n772_), .A2(new_n780_), .A3(new_n763_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n785_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n568_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n777_), .A2(new_n640_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n804_), .A2(new_n788_), .B1(new_n805_), .B2(new_n774_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n786_), .A2(KEYINPUT57), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n583_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n798_), .B(new_n799_), .C1(new_n808_), .C2(new_n793_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT118), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n795_), .A2(new_n811_), .A3(new_n798_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n804_), .A2(new_n788_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(new_n807_), .A3(new_n778_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n793_), .B1(new_n817_), .B2(new_n597_), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT117), .B(KEYINPUT59), .C1(new_n818_), .C2(new_n751_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n819_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n813_), .A2(KEYINPUT119), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT119), .B1(new_n813_), .B2(new_n820_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT120), .B(G113gat), .Z(new_n824_));
  NOR2_X1   g623(.A1(new_n460_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n797_), .B1(new_n823_), .B2(new_n825_), .ZN(G1340gat));
  INV_X1    g625(.A(G120gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n546_), .B2(KEYINPUT60), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n795_), .B(new_n828_), .C1(KEYINPUT60), .C2(new_n827_), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT121), .Z(new_n830_));
  AND3_X1   g629(.A1(new_n813_), .A2(new_n547_), .A3(new_n820_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n827_), .ZN(G1341gat));
  AOI21_X1  g631(.A(G127gat), .B1(new_n795_), .B2(new_n583_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n583_), .A2(KEYINPUT122), .A3(G127gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(KEYINPUT122), .B2(G127gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n823_), .B2(new_n835_), .ZN(G1342gat));
  AOI21_X1  g635(.A(G134gat), .B1(new_n795_), .B2(new_n594_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n640_), .A2(G134gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n823_), .B2(new_n838_), .ZN(G1343gat));
  NOR2_X1   g638(.A1(new_n818_), .A2(new_n616_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n589_), .A2(new_n623_), .A3(new_n308_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n459_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n547_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g646(.A1(new_n842_), .A2(KEYINPUT123), .A3(new_n597_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT123), .B1(new_n842_), .B2(new_n597_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT61), .B(G155gat), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1346gat));
  OAI21_X1  g652(.A(G162gat), .B1(new_n842_), .B2(new_n569_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n568_), .A2(G162gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n842_), .B2(new_n855_), .ZN(G1347gat));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n818_), .A2(new_n375_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n588_), .A2(new_n256_), .A3(new_n398_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n459_), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(G169gat), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n860_), .B2(G169gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n857_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n864_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(KEYINPUT62), .A3(new_n862_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n860_), .A2(new_n272_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(G1348gat));
  XOR2_X1   g668(.A(new_n858_), .B(KEYINPUT125), .Z(new_n870_));
  AND3_X1   g669(.A1(new_n859_), .A2(G176gat), .A3(new_n547_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n858_), .A2(new_n547_), .A3(new_n859_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n870_), .A2(new_n871_), .B1(new_n872_), .B2(new_n233_), .ZN(G1349gat));
  NAND2_X1  g672(.A1(new_n858_), .A2(new_n859_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n874_), .A2(new_n218_), .A3(new_n597_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n870_), .A2(new_n583_), .A3(new_n859_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n209_), .ZN(G1350gat));
  OAI21_X1  g676(.A(G190gat), .B1(new_n874_), .B2(new_n569_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n594_), .A2(new_n278_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n874_), .B2(new_n879_), .ZN(G1351gat));
  NOR3_X1   g679(.A1(new_n398_), .A2(new_n623_), .A3(new_n396_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n840_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n460_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT126), .B(G197gat), .Z(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1352gat));
  INV_X1    g684(.A(new_n882_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n547_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n583_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  AND2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n889_), .B2(new_n890_), .ZN(G1354gat));
  AOI21_X1  g692(.A(G218gat), .B1(new_n886_), .B2(new_n594_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n640_), .A2(G218gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT127), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n886_), .B2(new_n896_), .ZN(G1355gat));
endmodule


