//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_;
  INV_X1    g000(.A(G36gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G29gat), .ZN(new_n203_));
  INV_X1    g002(.A(G29gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G36gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G50gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G43gat), .ZN(new_n208_));
  INV_X1    g007(.A(G43gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G50gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n203_), .A2(new_n205_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(KEYINPUT15), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n213_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT73), .ZN(new_n218_));
  AND2_X1   g017(.A1(G1gat), .A2(G8gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT14), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G1gat), .A2(G8gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(KEYINPUT73), .A3(KEYINPUT14), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G1gat), .A2(G8gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT74), .B1(new_n219_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G1gat), .ZN(new_n228_));
  INV_X1    g027(.A(G8gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n222_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n225_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n225_), .A2(new_n233_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n214_), .B(new_n217_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n238_));
  AND4_X1   g037(.A1(new_n203_), .A2(new_n205_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n203_), .A2(new_n205_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G15gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G22gat), .ZN(new_n243_));
  INV_X1    g042(.A(G22gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G15gat), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n223_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n246_), .A2(new_n227_), .A3(new_n232_), .A4(new_n221_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n212_), .A2(KEYINPUT77), .A3(new_n213_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n241_), .A2(new_n247_), .A3(new_n248_), .A4(new_n234_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G229gat), .A2(G233gat), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n237_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n241_), .A2(new_n248_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(new_n236_), .B2(new_n235_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n250_), .B1(new_n253_), .B2(new_n249_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G113gat), .B(G141gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G169gat), .B(G197gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT78), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n255_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G78gat), .B(G106gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G22gat), .B(G50gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n262_), .B(new_n263_), .Z(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT3), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT2), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT87), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n271_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n272_), .A2(KEYINPUT1), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n272_), .B1(new_n273_), .B2(KEYINPUT1), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n276_), .B1(new_n277_), .B2(KEYINPUT86), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(KEYINPUT86), .B2(new_n277_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n266_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n268_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT29), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT88), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G197gat), .ZN(new_n286_));
  INV_X1    g085(.A(G204gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT89), .B(G197gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n288_), .B1(new_n289_), .B2(new_n287_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT90), .ZN(new_n292_));
  XOR2_X1   g091(.A(G211gat), .B(G218gat), .Z(new_n293_));
  INV_X1    g092(.A(KEYINPUT90), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n292_), .A2(KEYINPUT21), .A3(new_n293_), .A4(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n289_), .A2(new_n287_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT21), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n298_), .B1(G197gat), .B2(G204gat), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n293_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n291_), .B2(KEYINPUT21), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n296_), .A2(KEYINPUT91), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT91), .B1(new_n296_), .B2(new_n301_), .ZN(new_n304_));
  INV_X1    g103(.A(G228gat), .ZN(new_n305_));
  INV_X1    g104(.A(G233gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n303_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n282_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n285_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n296_), .A2(new_n301_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n283_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n275_), .A2(new_n315_), .A3(new_n281_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT28), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n314_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n265_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n310_), .A2(new_n314_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n317_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(new_n318_), .A3(new_n264_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT80), .ZN(new_n329_));
  INV_X1    g128(.A(G169gat), .ZN(new_n330_));
  INV_X1    g129(.A(G176gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(KEYINPUT24), .A3(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT25), .B(G183gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT79), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT26), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n335_), .B1(new_n336_), .B2(G190gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G190gat), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n334_), .B(new_n337_), .C1(new_n338_), .C2(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n333_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT81), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n342_), .A2(KEYINPUT23), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(KEYINPUT23), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(KEYINPUT24), .B2(new_n332_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n340_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT22), .B(G169gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n331_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n350_), .A2(new_n329_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n343_), .A2(KEYINPUT82), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n352_), .B(new_n344_), .Z(new_n353_));
  NOR2_X1   g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n351_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n348_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT30), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(new_n209_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT83), .B(G15gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n359_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G127gat), .B(G134gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G113gat), .B(G120gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT85), .B1(new_n368_), .B2(new_n369_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n373_), .B(KEYINPUT31), .Z(new_n374_));
  OR2_X1    g173(.A1(new_n357_), .A2(new_n358_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n375_), .A2(new_n359_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n367_), .B(new_n374_), .C1(new_n376_), .C2(new_n366_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n374_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n366_), .B1(new_n375_), .B2(new_n359_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n367_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G85gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT0), .B(G57gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n384_), .B(new_n385_), .Z(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n282_), .A2(new_n373_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n368_), .A2(new_n369_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n275_), .B(new_n281_), .C1(new_n371_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(KEYINPUT4), .A3(new_n390_), .ZN(new_n394_));
  XOR2_X1   g193(.A(KEYINPUT95), .B(KEYINPUT4), .Z(new_n395_));
  NAND3_X1  g194(.A1(new_n282_), .A2(new_n373_), .A3(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n387_), .B(new_n393_), .C1(new_n397_), .C2(new_n392_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n393_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n392_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n386_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n382_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT27), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n343_), .A2(new_n344_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n351_), .B1(new_n354_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n338_), .A2(new_n334_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n408_), .B(new_n409_), .C1(new_n332_), .C2(new_n407_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n406_), .B1(new_n353_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT20), .B1(new_n312_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n304_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n356_), .A2(new_n413_), .A3(new_n302_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT93), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n303_), .A2(new_n304_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT93), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n356_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n412_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT19), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n355_), .B(new_n348_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n312_), .B2(new_n411_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n421_), .ZN(new_n428_));
  XOR2_X1   g227(.A(G8gat), .B(G36gat), .Z(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G64gat), .B(G92gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n423_), .A2(new_n428_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n423_), .B2(new_n428_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n404_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT97), .B1(new_n427_), .B2(new_n421_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT97), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n424_), .A2(new_n439_), .A3(new_n422_), .A4(new_n426_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n438_), .B(new_n440_), .C1(new_n419_), .C2(new_n422_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n433_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n423_), .A2(new_n428_), .A3(new_n434_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(KEYINPUT27), .A3(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n437_), .A2(new_n444_), .A3(KEYINPUT98), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT98), .B1(new_n437_), .B2(new_n444_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n327_), .B(new_n403_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n402_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n448_), .A2(new_n437_), .A3(new_n444_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n423_), .A2(new_n428_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n433_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n394_), .A2(new_n392_), .A3(new_n396_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n387_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT33), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n401_), .ZN(new_n455_));
  OAI211_X1 g254(.A(KEYINPUT33), .B(new_n386_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n451_), .A2(new_n455_), .A3(new_n443_), .A4(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n434_), .A2(KEYINPUT32), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n441_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(KEYINPUT96), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n423_), .A2(new_n428_), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n402_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n326_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n382_), .B1(new_n449_), .B2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n261_), .B1(new_n447_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n471_));
  INV_X1    g270(.A(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G85gat), .ZN(new_n475_));
  INV_X1    g274(.A(G92gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT9), .A3(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(KEYINPUT9), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n470_), .A2(new_n474_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n478_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n482_), .B1(new_n486_), .B2(new_n470_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT8), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(new_n482_), .B2(KEYINPUT64), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n481_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n477_), .A2(new_n478_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n467_), .A2(new_n469_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n493_));
  INV_X1    g292(.A(G99gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n472_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n483_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n491_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT64), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT8), .B1(new_n491_), .B2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT65), .B1(new_n490_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n487_), .A2(new_n489_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n499_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT65), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .A4(new_n481_), .ZN(new_n505_));
  INV_X1    g304(.A(G64gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G57gat), .ZN(new_n507_));
  INV_X1    g306(.A(G57gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(G64gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n509_), .A3(KEYINPUT11), .ZN(new_n510_));
  INV_X1    g309(.A(G78gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(G71gat), .ZN(new_n512_));
  INV_X1    g311(.A(G71gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(G78gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G57gat), .B(G64gat), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n517_), .A2(KEYINPUT11), .A3(new_n512_), .A4(new_n514_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n501_), .A2(new_n505_), .A3(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(KEYINPUT12), .B(new_n520_), .C1(new_n516_), .C2(new_n518_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(new_n490_), .B2(new_n500_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n502_), .A2(new_n503_), .A3(new_n481_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT66), .B1(new_n528_), .B2(new_n524_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n522_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n501_), .A2(new_n505_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n521_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G230gat), .A2(G233gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n530_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n522_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n521_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n536_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G120gat), .B(G148gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(G176gat), .B(G204gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n542_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT13), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n547_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n525_), .A2(new_n526_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n528_), .A2(KEYINPUT66), .A3(new_n524_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n555_), .B(new_n522_), .C1(new_n539_), .C2(new_n531_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n540_), .B(new_n547_), .C1(new_n556_), .C2(new_n536_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(KEYINPUT13), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n550_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT69), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT76), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G127gat), .B(G155gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G183gat), .B(G211gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT17), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n235_), .A2(new_n236_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(new_n521_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(KEYINPUT17), .A3(new_n566_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT72), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n501_), .A2(new_n215_), .A3(new_n505_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT70), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n528_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .A4(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n581_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT35), .B1(new_n576_), .B2(new_n578_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n575_), .B(new_n583_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT71), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT36), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n587_), .A2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n576_), .A2(new_n578_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n584_), .B(new_n581_), .C1(new_n595_), .C2(KEYINPUT35), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n596_), .A2(new_n575_), .A3(new_n583_), .A4(new_n592_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n583_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(KEYINPUT36), .A3(new_n591_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT37), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n598_), .A2(new_n603_), .A3(new_n600_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  AND4_X1   g404(.A1(new_n465_), .A2(new_n560_), .A3(new_n574_), .A4(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n228_), .A3(new_n402_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n559_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n260_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n574_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT99), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n601_), .B1(new_n447_), .B2(new_n464_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n402_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n607_), .A2(new_n608_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n609_), .A2(new_n619_), .A3(new_n620_), .ZN(G1324gat));
  NOR2_X1   g420(.A1(new_n445_), .A2(new_n446_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n606_), .A2(new_n229_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n614_), .A2(new_n624_), .A3(new_n622_), .A4(new_n615_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(G8gat), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n614_), .A2(new_n622_), .A3(new_n615_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT100), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n626_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n627_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n623_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT40), .B(new_n623_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n617_), .B2(new_n382_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n638_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n382_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n606_), .A2(new_n242_), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n640_), .A3(new_n642_), .ZN(G1326gat));
  NAND2_X1  g442(.A1(new_n326_), .A2(new_n244_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT102), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n606_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n616_), .A2(new_n326_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(G22gat), .ZN(new_n649_));
  AOI211_X1 g448(.A(KEYINPUT42), .B(new_n244_), .C1(new_n616_), .C2(new_n326_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT103), .ZN(G1327gat));
  NAND2_X1  g451(.A1(new_n612_), .A2(new_n601_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n559_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n465_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n465_), .A2(KEYINPUT104), .A3(new_n654_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G29gat), .B1(new_n659_), .B2(new_n402_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n611_), .A2(new_n574_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n447_), .A2(new_n464_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n602_), .A2(new_n604_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT43), .B(new_n605_), .C1(new_n447_), .C2(new_n464_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT44), .B(new_n661_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n618_), .A2(new_n204_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n660_), .B1(new_n671_), .B2(new_n672_), .ZN(G1328gat));
  NAND4_X1  g472(.A1(new_n657_), .A2(new_n202_), .A3(new_n622_), .A4(new_n658_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT45), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n669_), .A2(new_n622_), .A3(new_n670_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G36gat), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT46), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n675_), .A2(new_n677_), .A3(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1329gat));
  NAND4_X1  g481(.A1(new_n669_), .A2(G43gat), .A3(new_n641_), .A4(new_n670_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n659_), .A2(new_n641_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(G43gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g485(.A1(new_n669_), .A2(new_n326_), .A3(new_n670_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G50gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n659_), .A2(new_n207_), .A3(new_n326_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT105), .ZN(G1331gat));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n663_), .B2(new_n261_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT106), .B(new_n260_), .C1(new_n447_), .C2(new_n464_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AND4_X1   g494(.A1(new_n559_), .A2(new_n695_), .A3(new_n574_), .A4(new_n605_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n508_), .A3(new_n402_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n560_), .A2(new_n260_), .A3(new_n612_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n615_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G57gat), .B1(new_n700_), .B2(new_n618_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n701_), .ZN(G1332gat));
  NAND3_X1  g501(.A1(new_n696_), .A2(new_n506_), .A3(new_n622_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n506_), .B1(new_n699_), .B2(new_n622_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT48), .Z(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1333gat));
  AOI21_X1  g505(.A(new_n513_), .B1(new_n699_), .B2(new_n641_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT49), .Z(new_n708_));
  NAND2_X1  g507(.A1(new_n641_), .A2(new_n513_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT107), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n696_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n708_), .A2(new_n711_), .ZN(G1334gat));
  NAND3_X1  g511(.A1(new_n696_), .A2(new_n511_), .A3(new_n326_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n511_), .B1(new_n699_), .B2(new_n326_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT50), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1335gat));
  NOR2_X1   g515(.A1(new_n560_), .A2(new_n653_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n695_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n475_), .A3(new_n402_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n665_), .A2(new_n666_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n610_), .A2(new_n260_), .A3(new_n574_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n402_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n720_), .B1(new_n725_), .B2(new_n475_), .ZN(G1336gat));
  NAND3_X1  g525(.A1(new_n719_), .A2(new_n476_), .A3(new_n622_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n622_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n729_), .B2(new_n476_), .ZN(G1337gat));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n641_), .B(new_n722_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G99gat), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n641_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n717_), .B(new_n734_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n731_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(KEYINPUT108), .A3(new_n735_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(KEYINPUT109), .A3(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n733_), .A2(new_n731_), .A3(new_n735_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n740_), .A2(new_n744_), .ZN(G1338gat));
  XNOR2_X1  g544(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n326_), .B(new_n722_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n749_), .B2(new_n472_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n327_), .A2(G106gat), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n717_), .B(new_n753_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n746_), .B1(new_n752_), .B2(new_n756_), .ZN(new_n757_));
  AND4_X1   g556(.A1(new_n756_), .A2(new_n751_), .A3(new_n750_), .A4(new_n746_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1339gat));
  INV_X1    g558(.A(G113gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n260_), .B2(KEYINPUT118), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n610_), .A2(new_n605_), .A3(new_n261_), .A4(new_n574_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT54), .Z(new_n763_));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n764_));
  INV_X1    g563(.A(new_n258_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n251_), .A2(new_n254_), .A3(new_n765_), .ZN(new_n766_));
  AND4_X1   g565(.A1(G229gat), .A2(new_n237_), .A3(G233gat), .A4(new_n249_), .ZN(new_n767_));
  AND4_X1   g566(.A1(new_n247_), .A2(new_n241_), .A3(new_n248_), .A4(new_n234_), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n248_), .A2(new_n241_), .B1(new_n247_), .B2(new_n234_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n250_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n765_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n767_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(KEYINPUT112), .A3(new_n765_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n766_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n557_), .A2(new_n764_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n764_), .B1(new_n557_), .B2(new_n775_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n536_), .B1(new_n530_), .B2(new_n534_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n537_), .B1(KEYINPUT55), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n556_), .A2(new_n781_), .A3(new_n536_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n551_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n501_), .A2(new_n505_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n786_), .A2(new_n521_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n532_), .A2(new_n533_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n531_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n790_), .A3(new_n535_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n535_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n781_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n537_), .A2(KEYINPUT55), .A3(new_n779_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(KEYINPUT56), .A3(new_n551_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n778_), .B1(new_n785_), .B2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT115), .B(new_n664_), .C1(new_n797_), .C2(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(KEYINPUT58), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n777_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n557_), .A2(new_n775_), .A3(new_n764_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n551_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n784_), .B(new_n547_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT115), .B1(new_n808_), .B2(new_n664_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT116), .B1(new_n800_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n601_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n260_), .A2(new_n557_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n785_), .B2(new_n796_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n548_), .A2(new_n775_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n811_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT57), .B(new_n811_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n817_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n664_), .B1(new_n797_), .B2(KEYINPUT58), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n799_), .A4(new_n798_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n815_), .A2(KEYINPUT113), .A3(new_n816_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n810_), .A2(new_n821_), .A3(new_n826_), .A4(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n763_), .B1(new_n828_), .B2(new_n612_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n622_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n830_), .A2(new_n402_), .A3(new_n327_), .A4(new_n641_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT59), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(KEYINPUT59), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n817_), .B1(new_n800_), .B2(new_n809_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n819_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT117), .B(new_n817_), .C1(new_n800_), .C2(new_n809_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n574_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n833_), .B1(new_n838_), .B2(new_n763_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n832_), .A2(new_n839_), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n761_), .B(new_n840_), .C1(KEYINPUT118), .C2(new_n760_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n828_), .A2(new_n612_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n763_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n831_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847_), .B2(new_n260_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n841_), .A2(new_n848_), .ZN(G1340gat));
  XOR2_X1   g648(.A(KEYINPUT119), .B(G120gat), .Z(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(KEYINPUT60), .B2(new_n850_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n846_), .A2(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT120), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n840_), .A2(new_n560_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n850_), .B2(new_n855_), .ZN(G1341gat));
  INV_X1    g655(.A(G127gat), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n574_), .B2(new_n858_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n859_), .B(new_n840_), .C1(new_n858_), .C2(new_n857_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G127gat), .B1(new_n847_), .B2(new_n574_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1342gat));
  NAND3_X1  g661(.A1(new_n832_), .A2(new_n839_), .A3(new_n664_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G134gat), .ZN(new_n864_));
  OR3_X1    g663(.A1(new_n846_), .A2(G134gat), .A3(new_n811_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n864_), .A2(new_n865_), .A3(KEYINPUT122), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1343gat));
  NOR3_X1   g669(.A1(new_n622_), .A2(new_n618_), .A3(new_n327_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n844_), .A2(new_n382_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n260_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g673(.A(new_n560_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g676(.A1(new_n829_), .A2(new_n641_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n871_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT123), .B1(new_n879_), .B2(new_n612_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n872_), .A2(new_n881_), .A3(new_n574_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n880_), .A2(new_n882_), .A3(new_n884_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1346gat));
  OR3_X1    g687(.A1(new_n879_), .A2(G162gat), .A3(new_n811_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G162gat), .B1(new_n879_), .B2(new_n605_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1347gat));
  NAND2_X1  g690(.A1(new_n834_), .A2(new_n835_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n818_), .A3(new_n837_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n763_), .B1(new_n893_), .B2(new_n612_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n622_), .A2(new_n403_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n326_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT125), .B1(new_n894_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n899_), .B(new_n896_), .C1(new_n838_), .C2(new_n763_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(new_n260_), .A3(new_n349_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n260_), .B(new_n896_), .C1(new_n838_), .C2(new_n763_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n330_), .B1(new_n905_), .B2(KEYINPUT124), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n903_), .B1(new_n906_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n894_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n910_), .A2(KEYINPUT124), .A3(new_n260_), .A4(new_n896_), .ZN(new_n911_));
  AND4_X1   g710(.A1(new_n903_), .A2(new_n911_), .A3(new_n908_), .A4(G169gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n902_), .B1(new_n909_), .B2(new_n912_), .ZN(G1348gat));
  NOR2_X1   g712(.A1(new_n829_), .A2(new_n326_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n895_), .A2(new_n331_), .A3(new_n560_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n901_), .A2(new_n559_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n917_), .A2(KEYINPUT126), .A3(new_n331_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n610_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(G176gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n916_), .B1(new_n918_), .B2(new_n921_), .ZN(G1349gat));
  NOR2_X1   g721(.A1(new_n895_), .A2(new_n612_), .ZN(new_n923_));
  AOI21_X1  g722(.A(G183gat), .B1(new_n914_), .B2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n612_), .A2(new_n334_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n901_), .B2(new_n925_), .ZN(G1350gat));
  INV_X1    g725(.A(new_n901_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G190gat), .B1(new_n927_), .B2(new_n605_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n901_), .A2(new_n338_), .A3(new_n601_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1351gat));
  NAND2_X1  g729(.A1(new_n622_), .A2(new_n448_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n878_), .A2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n261_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(new_n286_), .ZN(G1352gat));
  NOR2_X1   g734(.A1(new_n933_), .A2(new_n560_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(new_n287_), .ZN(G1353gat));
  NAND3_X1  g736(.A1(new_n878_), .A2(new_n574_), .A3(new_n932_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  AND2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n941_), .B1(new_n938_), .B2(new_n939_), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n933_), .B2(new_n605_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n811_), .A2(G218gat), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n878_), .A2(new_n932_), .A3(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(KEYINPUT127), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n943_), .A2(new_n948_), .A3(new_n945_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n949_), .ZN(G1355gat));
endmodule


