//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G57gat), .B(G64gat), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n203_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n202_), .B1(new_n205_), .B2(KEYINPUT11), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n213_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n219_), .A2(new_n220_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n214_), .B(KEYINPUT6), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT8), .B1(new_n227_), .B2(KEYINPUT64), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n214_), .ZN(new_n230_));
  OR2_X1    g029(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n231_));
  NAND2_X1  g030(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n231_), .A2(G99gat), .A3(G106gat), .A4(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n225_), .A2(new_n230_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n212_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n224_), .A2(new_n228_), .B1(new_n235_), .B2(KEYINPUT8), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n237_), .B(new_n226_), .C1(KEYINPUT9), .C2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT10), .B(G99gat), .Z(new_n240_));
  INV_X1    g039(.A(G106gat), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n211_), .B1(new_n236_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n209_), .A2(new_n210_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT8), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n225_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n212_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n247_), .B1(new_n234_), .B2(new_n212_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n245_), .B(new_n246_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n244_), .A2(new_n253_), .A3(KEYINPUT12), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n245_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT12), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n211_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n244_), .A2(new_n253_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(G230gat), .A3(G233gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n264_));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G176gat), .B(G204gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT66), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT68), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n260_), .A2(new_n262_), .A3(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT13), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT13), .B1(new_n272_), .B2(new_n273_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G232gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT34), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT35), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT70), .ZN(new_n284_));
  INV_X1    g083(.A(new_n282_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT35), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n236_), .A2(new_n243_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G43gat), .B(G50gat), .Z(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT71), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G43gat), .B(G50gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G29gat), .B(G36gat), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n290_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT15), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n290_), .A2(new_n293_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n294_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n290_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT15), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n287_), .B1(new_n288_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n302_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n255_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n284_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n295_), .A2(new_n296_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n288_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(KEYINPUT15), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n297_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n255_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n284_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n310_), .A2(new_n314_), .A3(new_n287_), .A4(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n308_), .A2(new_n316_), .A3(KEYINPUT72), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G190gat), .B(G218gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G134gat), .B(G162gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(KEYINPUT36), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n308_), .A2(new_n316_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(KEYINPUT36), .A3(new_n321_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n322_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n308_), .A2(new_n316_), .A3(KEYINPUT72), .A4(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n323_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT37), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n323_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT37), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G127gat), .B(G155gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(G211gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT16), .B(G183gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G231gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n246_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G15gat), .B(G22gat), .ZN(new_n340_));
  INV_X1    g139(.A(G1gat), .ZN(new_n341_));
  INV_X1    g140(.A(G8gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT14), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT73), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(new_n346_), .A3(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G1gat), .B(G8gat), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n339_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n337_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(KEYINPUT17), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n354_), .A2(new_n337_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT17), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n280_), .A2(new_n333_), .A3(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT19), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n368_));
  INV_X1    g167(.A(G204gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G197gat), .ZN(new_n370_));
  INV_X1    g169(.A(G197gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(G204gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT21), .ZN(new_n374_));
  OR2_X1    g173(.A1(G211gat), .A2(G218gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G211gat), .A2(G218gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G197gat), .B(G204gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT21), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n379_), .A2(new_n380_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT86), .B1(new_n373_), .B2(KEYINPUT21), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT86), .ZN(new_n383_));
  AOI211_X1 g182(.A(new_n383_), .B(new_n380_), .C1(new_n370_), .C2(new_n372_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n381_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(KEYINPUT87), .B(new_n381_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n378_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G183gat), .ZN(new_n397_));
  INV_X1    g196(.A(G183gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT25), .ZN(new_n399_));
  INV_X1    g198(.A(G190gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT26), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT26), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G190gat), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n397_), .A2(new_n399_), .A3(new_n401_), .A4(new_n403_), .ZN(new_n404_));
  OR3_X1    g203(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n405_));
  OR2_X1    g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(KEYINPUT24), .A3(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n395_), .A2(new_n404_), .A3(new_n405_), .A4(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G176gat), .ZN(new_n410_));
  AND2_X1   g209(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n413_), .B(new_n407_), .C1(new_n394_), .C2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n368_), .B1(new_n389_), .B2(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n401_), .A2(new_n403_), .ZN(new_n419_));
  OR3_X1    g218(.A1(new_n398_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n397_), .A2(KEYINPUT78), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n399_), .A4(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n405_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT79), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n408_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n408_), .A2(new_n424_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n422_), .B(new_n423_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n415_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n389_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n378_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n388_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n383_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n373_), .A2(KEYINPUT86), .A3(KEYINPUT21), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT87), .B1(new_n436_), .B2(new_n381_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n432_), .B1(new_n433_), .B2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT90), .B1(new_n438_), .B2(new_n428_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n367_), .B(new_n418_), .C1(new_n431_), .C2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT91), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n430_), .B1(new_n389_), .B2(new_n429_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(KEYINPUT90), .A3(new_n428_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n366_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(KEYINPUT91), .A3(new_n418_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n368_), .B1(new_n438_), .B2(new_n416_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n438_), .B2(new_n428_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n366_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n442_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G64gat), .B(G92gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(G8gat), .B(G36gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n442_), .A2(new_n446_), .A3(new_n455_), .A4(new_n449_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n364_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT98), .ZN(new_n460_));
  AOI221_X4 g259(.A(new_n378_), .B1(new_n416_), .B2(new_n460_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n417_), .A2(KEYINPUT98), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n443_), .A2(new_n444_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n464_));
  AOI21_X1  g263(.A(new_n367_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n448_), .A2(new_n366_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n456_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n467_), .A2(new_n458_), .A3(KEYINPUT27), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n459_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n428_), .B(KEYINPUT30), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT81), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G227gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT80), .ZN(new_n474_));
  XOR2_X1   g273(.A(G15gat), .B(G43gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(G71gat), .B(G99gat), .Z(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G127gat), .B(G134gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G113gat), .B(G120gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n480_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n486_), .B(KEYINPUT31), .Z(new_n487_));
  OR2_X1    g286(.A1(new_n470_), .A2(new_n471_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n488_), .A2(new_n472_), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n479_), .B(new_n487_), .C1(new_n489_), .C2(new_n478_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n487_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n478_), .B1(new_n488_), .B2(new_n472_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n479_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT99), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G225gat), .A2(G233gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT3), .ZN(new_n499_));
  INV_X1    g298(.A(G141gat), .ZN(new_n500_));
  INV_X1    g299(.A(G148gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G141gat), .A2(G148gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT2), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n502_), .A2(new_n505_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G155gat), .A2(G162gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(G155gat), .A2(G162gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n500_), .A2(new_n501_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(KEYINPUT1), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n510_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n509_), .A2(KEYINPUT1), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n512_), .B(new_n503_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n486_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n511_), .A2(new_n516_), .A3(new_n483_), .A4(new_n485_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  OR3_X1    g320(.A1(new_n517_), .A2(new_n486_), .A3(new_n519_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n498_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n518_), .A2(KEYINPUT4), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n522_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n524_), .B1(new_n525_), .B2(KEYINPUT4), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n523_), .B1(new_n526_), .B2(new_n498_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G1gat), .B(G29gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G85gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT0), .B(G57gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  OR2_X1    g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n498_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n523_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n496_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n532_), .A2(new_n496_), .A3(new_n535_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n495_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n517_), .A2(KEYINPUT29), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT82), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n540_), .B(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G22gat), .B(G50gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n517_), .A2(KEYINPUT29), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT85), .B1(new_n389_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(G233gat), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n550_), .A2(KEYINPUT84), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(KEYINPUT84), .ZN(new_n552_));
  OAI21_X1  g351(.A(G228gat), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT85), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n438_), .A2(new_n555_), .A3(new_n547_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n549_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n554_), .B1(new_n549_), .B2(new_n556_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT88), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G78gat), .B(G106gat), .Z(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n389_), .A2(KEYINPUT85), .A3(new_n548_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n555_), .B1(new_n438_), .B2(new_n547_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n553_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT88), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n549_), .A2(new_n556_), .A3(new_n554_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n559_), .A2(new_n561_), .A3(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n560_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT89), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n546_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n559_), .A2(new_n567_), .A3(KEYINPUT89), .A4(new_n561_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n564_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n571_), .A2(new_n572_), .B1(new_n574_), .B2(new_n546_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n469_), .A2(new_n539_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n538_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(new_n536_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n532_), .A2(new_n535_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n455_), .A2(KEYINPUT32), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n442_), .A2(new_n446_), .A3(new_n582_), .A4(new_n449_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n465_), .A2(new_n466_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n581_), .B(new_n583_), .C1(new_n584_), .C2(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n535_), .A2(KEYINPUT33), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT33), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n527_), .A2(new_n587_), .A3(new_n531_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n457_), .A2(new_n589_), .A3(new_n458_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n526_), .A2(new_n497_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT95), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT4), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n594_));
  NOR4_X1   g393(.A1(new_n594_), .A2(KEYINPUT95), .A3(new_n498_), .A4(new_n524_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n598_));
  INV_X1    g397(.A(new_n531_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n497_), .B1(new_n525_), .B2(KEYINPUT94), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(KEYINPUT94), .B2(new_n525_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .A4(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT95), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n526_), .B2(new_n497_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n599_), .B(new_n601_), .C1(new_n604_), .C2(new_n595_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT96), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n585_), .B1(new_n590_), .B2(new_n607_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n580_), .A2(new_n469_), .B1(new_n575_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n495_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n577_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n353_), .A2(new_n306_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n309_), .A2(new_n352_), .A3(new_n351_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n614_), .A2(KEYINPUT75), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT75), .B1(new_n614_), .B2(new_n615_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n613_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n612_), .B(KEYINPUT76), .Z(new_n619_));
  INV_X1    g418(.A(new_n353_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n615_), .B(new_n619_), .C1(new_n304_), .C2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT77), .B1(new_n618_), .B2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G169gat), .B(G197gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  AOI211_X1 g426(.A(KEYINPUT77), .B(new_n625_), .C1(new_n618_), .C2(new_n621_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n363_), .A2(new_n611_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n537_), .A2(new_n538_), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n630_), .A2(G1gat), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT101), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n362_), .A2(new_n331_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n276_), .A2(new_n277_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n629_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n611_), .A2(new_n636_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n341_), .B1(new_n641_), .B2(new_n579_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n632_), .B1(new_n633_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n635_), .A2(new_n643_), .ZN(G1324gat));
  OR2_X1    g443(.A1(new_n459_), .A2(new_n468_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n342_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n630_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n641_), .A2(KEYINPUT103), .A3(new_n645_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n640_), .B2(new_n469_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(G8gat), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n650_), .A2(KEYINPUT39), .A3(G8gat), .A4(new_n652_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n649_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  OAI21_X1  g458(.A(G15gat), .B1(new_n640_), .B2(new_n495_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT41), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n630_), .A2(G15gat), .A3(new_n495_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n640_), .B2(new_n575_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n575_), .A2(G22gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n630_), .B2(new_n666_), .ZN(G1327gat));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n568_), .A2(new_n570_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n545_), .A3(new_n572_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n574_), .A2(new_n546_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n469_), .A2(new_n672_), .A3(new_n631_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n608_), .A2(new_n575_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n576_), .B1(new_n675_), .B2(new_n495_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n331_), .B(new_n329_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n668_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n610_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT43), .B(new_n333_), .C1(new_n679_), .C2(new_n576_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n678_), .A2(new_n362_), .A3(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT106), .B1(KEYINPUT105), .B2(KEYINPUT44), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(KEYINPUT106), .B2(KEYINPUT44), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n681_), .A2(new_n639_), .A3(new_n683_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n678_), .A2(new_n362_), .A3(new_n639_), .A4(new_n680_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n682_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n684_), .A2(new_n579_), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G29gat), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n676_), .A2(new_n638_), .A3(new_n637_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n361_), .A2(new_n328_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(G29gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n631_), .B2(new_n692_), .ZN(G1328gat));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n645_), .A3(new_n686_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  INV_X1    g494(.A(G36gat), .ZN(new_n696_));
  AND4_X1   g495(.A1(new_n696_), .A2(new_n689_), .A3(new_n645_), .A4(new_n690_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n695_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n695_), .A2(new_n699_), .A3(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  NAND4_X1  g503(.A1(new_n684_), .A2(G43gat), .A3(new_n610_), .A4(new_n686_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n691_), .A2(new_n495_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(G43gat), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g507(.A1(new_n691_), .A2(G50gat), .A3(new_n575_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n684_), .A2(new_n672_), .A3(new_n686_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(G50gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G50gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(G1331gat));
  NAND4_X1  g513(.A1(new_n611_), .A2(new_n638_), .A3(new_n280_), .A4(new_n636_), .ZN(new_n715_));
  INV_X1    g514(.A(G57gat), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n631_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n333_), .A2(new_n278_), .A3(new_n362_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n718_), .A2(KEYINPUT109), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(KEYINPUT109), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n719_), .A2(new_n611_), .A3(new_n638_), .A4(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT110), .Z(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n579_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n717_), .B1(new_n723_), .B2(new_n716_), .ZN(G1332gat));
  OAI21_X1  g523(.A(G64gat), .B1(new_n715_), .B2(new_n469_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT48), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n469_), .A2(G64gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n721_), .B2(new_n727_), .ZN(G1333gat));
  OAI21_X1  g527(.A(G71gat), .B1(new_n715_), .B2(new_n495_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT111), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(KEYINPUT111), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n732_), .A2(KEYINPUT49), .ZN(new_n733_));
  OR3_X1    g532(.A1(new_n721_), .A2(G71gat), .A3(new_n495_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n730_), .A2(KEYINPUT49), .A3(new_n731_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(G1334gat));
  OAI21_X1  g535(.A(G78gat), .B1(new_n715_), .B2(new_n575_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT50), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n575_), .A2(G78gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n721_), .B2(new_n739_), .ZN(G1335gat));
  NAND3_X1  g539(.A1(new_n681_), .A2(new_n638_), .A3(new_n637_), .ZN(new_n741_));
  INV_X1    g540(.A(G85gat), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n631_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n611_), .A2(new_n638_), .A3(new_n280_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n746_), .B2(new_n690_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n690_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n745_), .A2(KEYINPUT112), .A3(new_n748_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n579_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n743_), .B1(new_n751_), .B2(new_n742_), .ZN(G1336gat));
  AOI21_X1  g551(.A(G92gat), .B1(new_n750_), .B2(new_n645_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n741_), .A2(new_n469_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(G92gat), .B2(new_n754_), .ZN(G1337gat));
  OAI21_X1  g554(.A(G99gat), .B1(new_n741_), .B2(new_n495_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n610_), .B(new_n240_), .C1(new_n747_), .C2(new_n749_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n759_), .A2(KEYINPUT51), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(KEYINPUT51), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n758_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n756_), .A2(new_n757_), .A3(new_n759_), .A4(KEYINPUT51), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1338gat));
  OAI211_X1 g563(.A(new_n241_), .B(new_n672_), .C1(new_n747_), .C2(new_n749_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n678_), .A2(new_n638_), .A3(new_n362_), .A4(new_n680_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n766_), .A2(new_n575_), .A3(new_n278_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n767_), .A2(KEYINPUT52), .A3(new_n241_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n681_), .A2(new_n672_), .A3(new_n638_), .A4(new_n637_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n765_), .B1(new_n768_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n765_), .C1(new_n768_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  NOR4_X1   g575(.A1(new_n645_), .A2(new_n672_), .A3(new_n631_), .A4(new_n495_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n263_), .A2(new_n268_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(KEYINPUT114), .A2(G230gat), .A3(G233gat), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(new_n780_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n781_), .B1(new_n260_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n258_), .A2(KEYINPUT55), .A3(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n268_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n786_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n258_), .A2(KEYINPUT55), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n254_), .A2(new_n257_), .B1(G230gat), .B2(G233gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n784_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n268_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n629_), .B(new_n779_), .C1(new_n790_), .C2(new_n796_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n618_), .A2(new_n621_), .A3(new_n626_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n614_), .A2(new_n615_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT75), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n614_), .A2(new_n615_), .A3(KEYINPUT75), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n619_), .A3(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n615_), .B1(new_n304_), .B2(new_n620_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n619_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n626_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT115), .B1(new_n798_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n806_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n625_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n618_), .A2(new_n621_), .A3(new_n626_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n808_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n274_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n797_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT57), .B1(new_n816_), .B2(new_n328_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n818_), .B(new_n331_), .C1(new_n797_), .C2(new_n815_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n789_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n795_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n778_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT58), .B1(new_n823_), .B2(new_n814_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT116), .B1(new_n824_), .B2(new_n677_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n814_), .B(new_n779_), .C1(new_n790_), .C2(new_n796_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n333_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n823_), .A2(KEYINPUT58), .A3(new_n814_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n825_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n361_), .B1(new_n820_), .B2(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n330_), .A2(new_n361_), .A3(new_n638_), .A4(new_n332_), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n834_), .A2(new_n637_), .A3(KEYINPUT54), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT54), .B1(new_n834_), .B2(new_n637_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n777_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G113gat), .B1(new_n839_), .B2(new_n629_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n838_), .A2(KEYINPUT117), .A3(KEYINPUT59), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT117), .B1(new_n838_), .B2(KEYINPUT59), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT59), .B1(new_n777_), .B2(KEYINPUT118), .ZN(new_n844_));
  OAI221_X1 g643(.A(new_n844_), .B1(KEYINPUT118), .B2(new_n777_), .C1(new_n833_), .C2(new_n837_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n843_), .A2(G113gat), .A3(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n840_), .B1(new_n846_), .B2(new_n629_), .ZN(G1340gat));
  NAND4_X1  g646(.A1(new_n843_), .A2(KEYINPUT121), .A3(new_n280_), .A4(new_n845_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n838_), .A2(KEYINPUT59), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n838_), .A2(KEYINPUT117), .A3(KEYINPUT59), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n851_), .A2(new_n280_), .A3(new_n845_), .A4(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT119), .B(G120gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n848_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT60), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n856_), .B1(new_n637_), .B2(new_n858_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT120), .Z(new_n861_));
  NAND3_X1  g660(.A1(new_n839_), .A2(new_n859_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n862_), .ZN(G1341gat));
  AOI21_X1  g662(.A(G127gat), .B1(new_n839_), .B2(new_n361_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n843_), .A2(G127gat), .A3(new_n845_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n361_), .ZN(G1342gat));
  AOI21_X1  g665(.A(G134gat), .B1(new_n839_), .B2(new_n331_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n843_), .A2(new_n333_), .A3(new_n845_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g668(.A1(new_n820_), .A2(new_n832_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n362_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n835_), .A2(new_n836_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n610_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n579_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n645_), .A2(new_n575_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n629_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n280_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n361_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  AOI21_X1  g683(.A(G162gat), .B1(new_n877_), .B2(new_n331_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n874_), .A2(new_n677_), .A3(new_n876_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(G162gat), .B2(new_n886_), .ZN(G1347gat));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n469_), .A2(new_n672_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n539_), .B(new_n889_), .C1(new_n833_), .C2(new_n837_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n629_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n888_), .B1(new_n892_), .B2(G169gat), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n888_), .B(G169gat), .C1(new_n890_), .C2(new_n638_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(KEYINPUT62), .A3(new_n895_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n891_), .B(new_n629_), .C1(new_n412_), .C2(new_n411_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n893_), .B2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n896_), .A2(new_n897_), .A3(new_n900_), .ZN(G1348gat));
  OAI21_X1  g700(.A(new_n410_), .B1(new_n890_), .B2(new_n278_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n890_), .A2(new_n410_), .ZN(new_n903_));
  AOI21_X1  g702(.A(KEYINPUT123), .B1(new_n903_), .B2(new_n280_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905_));
  INV_X1    g704(.A(new_n280_), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n890_), .A2(new_n905_), .A3(new_n410_), .A4(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n902_), .B1(new_n904_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT124), .B(new_n902_), .C1(new_n904_), .C2(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1349gat));
  NOR2_X1   g711(.A1(new_n890_), .A2(new_n362_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n398_), .A2(KEYINPUT125), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n913_), .A2(new_n397_), .A3(new_n399_), .A4(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(KEYINPUT125), .A2(G183gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n913_), .B2(new_n916_), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n890_), .B2(new_n677_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n331_), .A2(new_n419_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n890_), .B2(new_n919_), .ZN(G1351gat));
  NAND2_X1  g719(.A1(new_n873_), .A2(new_n580_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n921_), .A2(new_n469_), .A3(new_n638_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT126), .B(G197gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1352gat));
  NOR3_X1   g723(.A1(new_n921_), .A2(new_n469_), .A3(new_n906_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1353gat));
  INV_X1    g726(.A(new_n921_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n928_), .A2(new_n645_), .A3(new_n361_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT63), .B(G211gat), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n929_), .B2(new_n932_), .ZN(G1354gat));
  INV_X1    g732(.A(G218gat), .ZN(new_n934_));
  NOR4_X1   g733(.A1(new_n921_), .A2(new_n934_), .A3(new_n469_), .A4(new_n677_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n928_), .A2(new_n645_), .A3(new_n331_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n934_), .B2(new_n936_), .ZN(G1355gat));
endmodule


