//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT89), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n205_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(new_n203_), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n207_), .B(new_n209_), .Z(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  OR2_X1    g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT22), .B(G169gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT91), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n211_), .B(new_n215_), .C1(new_n217_), .C2(G176gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n219_), .B1(new_n212_), .B2(KEYINPUT23), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n212_), .A2(KEYINPUT23), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n211_), .A2(KEYINPUT24), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  MUX2_X1   g023(.A(new_n223_), .B(KEYINPUT24), .S(new_n224_), .Z(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT25), .B(G183gat), .Z(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT26), .B(G190gat), .Z(new_n227_));
  OAI211_X1 g026(.A(new_n222_), .B(new_n225_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n210_), .A2(new_n218_), .A3(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n229_), .A2(KEYINPUT20), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT92), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G226gat), .A2(G233gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT19), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n210_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n226_), .A2(new_n227_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(KEYINPUT77), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(KEYINPUT77), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n237_), .A2(new_n213_), .A3(new_n238_), .A4(new_n225_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n222_), .A2(new_n214_), .ZN(new_n240_));
  INV_X1    g039(.A(G169gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT79), .B1(new_n241_), .B2(KEYINPUT22), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT78), .B(KEYINPUT22), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n243_), .B2(G169gat), .ZN(new_n244_));
  INV_X1    g043(.A(G176gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(G169gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n245_), .B1(new_n246_), .B2(KEYINPUT79), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n240_), .B(new_n211_), .C1(new_n244_), .C2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n239_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n235_), .A2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n230_), .A2(new_n231_), .A3(new_n234_), .A4(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n250_), .A2(KEYINPUT20), .A3(new_n234_), .A4(new_n229_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT92), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G8gat), .B(G36gat), .Z(new_n255_));
  XNOR2_X1  g054(.A(G64gat), .B(G92gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT20), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n218_), .A2(new_n228_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n235_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n210_), .A2(new_n248_), .A3(new_n239_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n233_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n254_), .A2(new_n260_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n260_), .B1(new_n254_), .B2(new_n266_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n202_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G1gat), .B(G29gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(G57gat), .B(G85gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  XOR2_X1   g074(.A(G127gat), .B(G134gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT84), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G113gat), .B(G120gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT88), .ZN(new_n283_));
  INV_X1    g082(.A(G141gat), .ZN(new_n284_));
  INV_X1    g083(.A(G148gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR3_X1   g085(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n288_));
  AOI22_X1  g087(.A1(KEYINPUT2), .A2(new_n286_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n283_), .B(new_n289_), .C1(new_n288_), .C2(new_n287_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n291_), .B(KEYINPUT86), .Z(new_n292_));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n293_), .B(KEYINPUT1), .Z(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n286_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n284_), .A2(new_n285_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n280_), .A2(new_n281_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G225gat), .A2(G233gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n300_), .A2(KEYINPUT94), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n305_), .A2(new_n279_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n279_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n304_), .B1(new_n308_), .B2(KEYINPUT4), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n305_), .B(new_n280_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(new_n303_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n275_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n302_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n275_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n310_), .A2(new_n281_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n313_), .B(new_n314_), .C1(new_n315_), .C2(new_n304_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n233_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n230_), .A2(new_n250_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n320_), .B2(new_n233_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n202_), .B1(new_n321_), .B2(new_n259_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT96), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n267_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n322_), .B2(new_n267_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n270_), .B(new_n318_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT85), .ZN(new_n328_));
  XOR2_X1   g127(.A(G15gat), .B(G43gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT82), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G71gat), .B(G99gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G227gat), .A2(G233gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n333_), .B(KEYINPUT83), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n332_), .B(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n336_));
  NAND2_X1  g135(.A1(new_n249_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n249_), .A2(new_n336_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n335_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n335_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n328_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n334_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n332_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n339_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n337_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n340_), .A2(new_n347_), .A3(KEYINPUT85), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n279_), .B(KEYINPUT31), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n343_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n349_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n328_), .B(new_n351_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n300_), .A2(KEYINPUT29), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G228gat), .A2(G233gat), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n354_), .A2(new_n235_), .B1(KEYINPUT90), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT90), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n354_), .A2(new_n235_), .A3(new_n358_), .A4(new_n357_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G78gat), .B(G106gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G22gat), .B(G50gat), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n360_), .A2(new_n361_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n362_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n366_), .B1(new_n371_), .B2(new_n363_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n300_), .A2(KEYINPUT29), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT28), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n368_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n374_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n367_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n371_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n353_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n374_), .B1(new_n368_), .B2(new_n372_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n350_), .A2(new_n352_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(new_n378_), .A3(new_n376_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n321_), .A2(KEYINPUT32), .A3(new_n260_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n260_), .A2(KEYINPUT32), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n254_), .A2(new_n266_), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n317_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT33), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n316_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n309_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n392_), .A2(KEYINPUT33), .A3(new_n313_), .A4(new_n314_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n301_), .A2(new_n302_), .ZN(new_n394_));
  OAI221_X1 g193(.A(new_n275_), .B1(new_n310_), .B2(new_n302_), .C1(new_n315_), .C2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n268_), .A2(new_n269_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n389_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n353_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n327_), .A2(new_n385_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G120gat), .B(G148gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT5), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G176gat), .B(G204gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G85gat), .A2(G92gat), .ZN(new_n406_));
  AND2_X1   g205(.A1(G85gat), .A2(G92gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(KEYINPUT9), .ZN(new_n408_));
  INV_X1    g207(.A(G92gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT67), .ZN(new_n410_));
  INV_X1    g209(.A(G85gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(KEYINPUT67), .A2(G85gat), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n409_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT9), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT66), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT66), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT9), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n408_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT68), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT68), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n422_), .B(new_n408_), .C1(new_n414_), .C2(new_n419_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G99gat), .A2(G106gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n426_));
  NOR2_X1   g225(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n429_));
  NAND2_X1  g228(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n424_), .A3(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT65), .B(G106gat), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n428_), .A2(new_n431_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n421_), .A2(new_n423_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT8), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n428_), .A2(new_n431_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G99gat), .A2(G106gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(KEYINPUT70), .A2(KEYINPUT7), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  OAI22_X1  g242(.A1(KEYINPUT70), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n440_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n407_), .A2(new_n406_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n439_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  AOI211_X1 g248(.A(KEYINPUT8), .B(new_n449_), .C1(new_n440_), .C2(new_n445_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n437_), .B(new_n438_), .C1(new_n448_), .C2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G57gat), .B(G64gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT11), .ZN(new_n453_));
  XOR2_X1   g252(.A(G71gat), .B(G78gat), .Z(new_n454_));
  OR2_X1    g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n452_), .A2(KEYINPUT11), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n454_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n455_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n443_), .A2(new_n444_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT8), .B1(new_n461_), .B2(new_n449_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n446_), .A2(new_n439_), .A3(new_n447_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n423_), .A2(new_n436_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n462_), .A2(new_n463_), .B1(new_n464_), .B2(new_n421_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT71), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT12), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n451_), .B(new_n459_), .C1(new_n465_), .C2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n437_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n469_), .A2(new_n466_), .A3(KEYINPUT12), .A4(new_n458_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G230gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT64), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n465_), .A2(new_n458_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n469_), .A2(new_n459_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n474_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n405_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n473_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n481_), .A2(new_n478_), .A3(new_n404_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT13), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT13), .B1(new_n480_), .B2(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G113gat), .B(G141gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT76), .ZN(new_n490_));
  XOR2_X1   g289(.A(G169gat), .B(G197gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT74), .B(G8gat), .Z(new_n493_));
  INV_X1    g292(.A(G1gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT14), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT73), .B(G15gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G22gat), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n496_), .A2(G22gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G1gat), .B(G8gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n495_), .A2(new_n498_), .A3(new_n497_), .A4(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G29gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G229gat), .A2(G233gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n507_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n502_), .A2(new_n511_), .A3(new_n503_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n508_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(KEYINPUT15), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT15), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n507_), .A2(new_n516_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n515_), .A2(new_n502_), .A3(new_n517_), .A4(new_n503_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n510_), .B1(new_n508_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n492_), .B1(new_n514_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n492_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n513_), .A3(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n488_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n400_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n458_), .B(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n529_), .B(new_n504_), .Z(new_n530_));
  XNOR2_X1  g329(.A(G127gat), .B(G155gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT16), .ZN(new_n532_));
  XOR2_X1   g331(.A(G183gat), .B(G211gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n534_), .A2(KEYINPUT71), .A3(new_n535_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT75), .ZN(new_n540_));
  INV_X1    g339(.A(new_n538_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n537_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT34), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n469_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n552_));
  OAI22_X1  g351(.A1(new_n469_), .A2(new_n511_), .B1(KEYINPUT35), .B2(new_n548_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n465_), .A2(new_n507_), .B1(new_n550_), .B2(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n551_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n469_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT36), .Z(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(KEYINPUT36), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n554_), .A2(new_n558_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n566_), .B2(KEYINPUT72), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n564_), .B(new_n566_), .C1(KEYINPUT72), .C2(new_n568_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n546_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n527_), .A2(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT97), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(KEYINPUT97), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(new_n494_), .A3(new_n317_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT38), .ZN(new_n579_));
  INV_X1    g378(.A(new_n567_), .ZN(new_n580_));
  NOR4_X1   g379(.A1(new_n400_), .A2(new_n580_), .A3(new_n526_), .A4(new_n539_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n581_), .A2(new_n317_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n579_), .B1(new_n494_), .B2(new_n582_), .ZN(G1324gat));
  OAI21_X1  g382(.A(new_n270_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT99), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT99), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(G8gat), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n575_), .A2(new_n584_), .A3(new_n493_), .A4(new_n576_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n592_), .A2(KEYINPUT98), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(KEYINPUT98), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n590_), .B(new_n591_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(G1325gat));
  INV_X1    g396(.A(G15gat), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n577_), .A2(new_n598_), .A3(new_n353_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n581_), .B2(new_n353_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(G1326gat));
  INV_X1    g402(.A(G22gat), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n375_), .A2(new_n379_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n581_), .B2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT42), .Z(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n604_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT102), .Z(new_n609_));
  NAND2_X1  g408(.A1(new_n577_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(G1327gat));
  XNOR2_X1  g410(.A(new_n572_), .B(KEYINPUT103), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT43), .B1(new_n400_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n398_), .A2(new_n399_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n382_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n614_), .B1(new_n617_), .B2(new_n326_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT43), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(new_n572_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n545_), .B1(new_n613_), .B2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(KEYINPUT44), .A3(new_n525_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(G29gat), .A3(new_n317_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT44), .B1(new_n621_), .B2(new_n525_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n545_), .A2(new_n567_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n527_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(new_n318_), .ZN(new_n627_));
  OAI22_X1  g426(.A1(new_n623_), .A2(new_n624_), .B1(G29gat), .B2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT104), .Z(G1328gat));
  INV_X1    g428(.A(KEYINPUT106), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT46), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT107), .ZN(new_n634_));
  INV_X1    g433(.A(new_n612_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n619_), .B1(new_n618_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n572_), .A2(new_n619_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n400_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n525_), .B(new_n546_), .C1(new_n636_), .C2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n584_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G36gat), .B1(new_n641_), .B2(new_n624_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT105), .B(G36gat), .C1(new_n641_), .C2(new_n624_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n584_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(G36gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n527_), .A2(new_n625_), .A3(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT45), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n630_), .A2(new_n631_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n634_), .B1(new_n646_), .B2(new_n653_), .ZN(new_n654_));
  AOI211_X1 g453(.A(KEYINPUT107), .B(new_n652_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n633_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n645_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n639_), .A2(new_n640_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n622_), .A3(new_n584_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT105), .B1(new_n659_), .B2(G36gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n653_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT107), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n646_), .A2(new_n634_), .A3(new_n653_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n632_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n656_), .A2(new_n664_), .ZN(G1329gat));
  AND2_X1   g464(.A1(new_n658_), .A2(new_n622_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(G43gat), .A3(new_n353_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n626_), .A2(new_n382_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(G43gat), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g469(.A(new_n666_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n605_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G50gat), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(G50gat), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT108), .Z(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n626_), .B2(new_n675_), .ZN(G1331gat));
  NAND2_X1  g475(.A1(new_n573_), .A2(new_n488_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n524_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n400_), .B(new_n679_), .C1(new_n678_), .C2(new_n677_), .ZN(new_n680_));
  INV_X1    g479(.A(G57gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(new_n681_), .A3(new_n317_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n540_), .A2(new_n544_), .A3(new_n524_), .ZN(new_n683_));
  OR4_X1    g482(.A1(new_n580_), .A2(new_n400_), .A3(new_n487_), .A4(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n318_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(G1332gat));
  OAI21_X1  g485(.A(G64gat), .B1(new_n684_), .B2(new_n647_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n647_), .A2(G64gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT111), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n680_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(G1333gat));
  OAI21_X1  g492(.A(G71gat), .B1(new_n684_), .B2(new_n382_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT49), .ZN(new_n695_));
  INV_X1    g494(.A(G71gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n680_), .A2(new_n696_), .A3(new_n353_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1334gat));
  OAI21_X1  g497(.A(G78gat), .B1(new_n684_), .B2(new_n672_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT50), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n672_), .A2(G78gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT112), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n680_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(G1335gat));
  NAND2_X1  g503(.A1(new_n520_), .A2(new_n523_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n487_), .A2(new_n705_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n618_), .A2(new_n625_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G85gat), .B1(new_n707_), .B2(new_n317_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n621_), .A2(new_n706_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n318_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n710_), .B2(new_n711_), .ZN(G1336gat));
  OAI21_X1  g511(.A(G92gat), .B1(new_n709_), .B2(new_n647_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n707_), .A2(new_n409_), .A3(new_n584_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1337gat));
  NOR2_X1   g514(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n716_));
  OAI21_X1  g515(.A(G99gat), .B1(new_n709_), .B2(new_n382_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n707_), .A2(new_n434_), .A3(new_n353_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n719_), .B(new_n720_), .Z(G1338gat));
  OAI21_X1  g520(.A(G106gat), .B1(new_n709_), .B2(new_n672_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT52), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n707_), .A2(new_n435_), .A3(new_n605_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g525(.A1(new_n647_), .A2(new_n317_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n380_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT121), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT117), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT57), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n508_), .A2(new_n512_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n492_), .B1(new_n733_), .B2(new_n509_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n508_), .A2(new_n510_), .A3(new_n518_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n520_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n483_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n475_), .A2(new_n479_), .A3(new_n405_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT116), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n705_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n740_), .B2(new_n705_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n468_), .A2(new_n473_), .A3(new_n470_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n481_), .B2(KEYINPUT55), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n748_), .B(new_n473_), .C1(new_n468_), .C2(new_n470_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n404_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT56), .B(new_n404_), .C1(new_n747_), .C2(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n739_), .B1(new_n745_), .B2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n731_), .B(new_n732_), .C1(new_n755_), .C2(new_n580_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n731_), .A2(new_n732_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT116), .B1(new_n524_), .B2(new_n482_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n742_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n567_), .B(new_n757_), .C1(new_n760_), .C2(new_n739_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n756_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n737_), .A2(new_n740_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n475_), .A2(new_n748_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n481_), .A2(KEYINPUT55), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n746_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n404_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n753_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT58), .B(new_n764_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT119), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n763_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT119), .A3(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT118), .B(new_n572_), .C1(new_n773_), .C2(KEYINPUT58), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n572_), .B1(new_n773_), .B2(KEYINPUT58), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT118), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n775_), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT120), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n762_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AND4_X1   g581(.A1(KEYINPUT119), .A2(new_n754_), .A3(KEYINPUT58), .A4(new_n764_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT119), .B1(new_n773_), .B2(KEYINPUT58), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n764_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT118), .B1(new_n788_), .B2(new_n572_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n776_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n785_), .B(new_n781_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n730_), .B1(new_n782_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n785_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT120), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n795_), .A2(KEYINPUT121), .A3(new_n791_), .A4(new_n762_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n539_), .A3(new_n796_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n683_), .A2(KEYINPUT114), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n683_), .A2(KEYINPUT114), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801_));
  INV_X1    g600(.A(new_n572_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n487_), .A4(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n488_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n806_), .A2(KEYINPUT115), .A3(new_n801_), .A4(new_n802_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n800_), .A2(new_n487_), .A3(new_n802_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT54), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(new_n807_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n729_), .B1(new_n797_), .B2(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n811_), .A2(KEYINPUT122), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(KEYINPUT122), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(G113gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n705_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n805_), .A2(new_n807_), .A3(new_n809_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n545_), .B1(new_n762_), .B2(new_n794_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n729_), .A2(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n811_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(G113gat), .B1(new_n823_), .B2(new_n524_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n816_), .A2(new_n824_), .ZN(G1340gat));
  INV_X1    g624(.A(KEYINPUT60), .ZN(new_n826_));
  INV_X1    g625(.A(G120gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n488_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n814_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(G120gat), .B1(new_n823_), .B2(new_n487_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1341gat));
  INV_X1    g631(.A(G127gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n814_), .A2(new_n833_), .A3(new_n545_), .ZN(new_n834_));
  OAI21_X1  g633(.A(G127gat), .B1(new_n823_), .B2(new_n539_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1342gat));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n837_));
  NOR4_X1   g636(.A1(new_n812_), .A2(new_n813_), .A3(G134gat), .A4(new_n567_), .ZN(new_n838_));
  INV_X1    g637(.A(G134gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n796_), .A2(new_n539_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n756_), .A2(new_n761_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n794_), .B2(KEYINPUT120), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT121), .B1(new_n842_), .B2(new_n791_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n810_), .B1(new_n840_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n728_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n845_), .A2(KEYINPUT59), .B1(new_n819_), .B2(new_n820_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n839_), .B1(new_n846_), .B2(new_n572_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n837_), .B1(new_n838_), .B2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n814_), .A2(new_n839_), .A3(new_n580_), .ZN(new_n849_));
  OAI21_X1  g648(.A(G134gat), .B1(new_n823_), .B2(new_n802_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n850_), .A3(KEYINPUT123), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(G1343gat));
  AOI21_X1  g651(.A(new_n384_), .B1(new_n797_), .B2(new_n810_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n727_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n705_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n488_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n844_), .A2(new_n615_), .A3(new_n545_), .A4(new_n854_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n853_), .A2(KEYINPUT124), .A3(new_n545_), .A4(new_n854_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n860_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n863_), .A2(new_n865_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT125), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n863_), .A2(new_n865_), .A3(new_n864_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n860_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n868_), .A2(new_n873_), .ZN(G1346gat));
  AOI21_X1  g673(.A(G162gat), .B1(new_n855_), .B2(new_n580_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n635_), .A2(G162gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n855_), .B2(new_n876_), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n647_), .A2(new_n317_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n353_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n605_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G169gat), .B1(new_n881_), .B2(new_n524_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n882_), .A2(KEYINPUT62), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(KEYINPUT62), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n881_), .B(KEYINPUT126), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n524_), .A2(new_n217_), .ZN(new_n886_));
  OAI22_X1  g685(.A1(new_n883_), .A2(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(G1348gat));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n881_), .B(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G176gat), .B1(new_n889_), .B2(new_n488_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n844_), .A2(new_n672_), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n891_), .A2(new_n245_), .A3(new_n487_), .A4(new_n879_), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT127), .B1(new_n890_), .B2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n245_), .B1(new_n885_), .B2(new_n487_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n892_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n893_), .A2(new_n897_), .ZN(G1349gat));
  OR3_X1    g697(.A1(new_n891_), .A2(new_n546_), .A3(new_n879_), .ZN(new_n899_));
  INV_X1    g698(.A(G183gat), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n542_), .A2(new_n226_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n899_), .A2(new_n900_), .B1(new_n889_), .B2(new_n901_), .ZN(G1350gat));
  OAI21_X1  g701(.A(G190gat), .B1(new_n885_), .B2(new_n802_), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n567_), .A2(new_n227_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n885_), .B2(new_n904_), .ZN(G1351gat));
  NAND2_X1  g704(.A1(new_n853_), .A2(new_n878_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n705_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n488_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g710(.A1(new_n906_), .A2(new_n539_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  AND2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n915_), .B1(new_n912_), .B2(new_n913_), .ZN(G1354gat));
  OAI21_X1  g715(.A(G218gat), .B1(new_n906_), .B2(new_n802_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n567_), .A2(G218gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n906_), .B2(new_n918_), .ZN(G1355gat));
endmodule


