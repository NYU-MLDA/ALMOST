//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  XOR2_X1   g001(.A(G120gat), .B(G148gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G176gat), .B(G204gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT8), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT7), .ZN(new_n209_));
  INV_X1    g008(.A(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(KEYINPUT6), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT6), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT65), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n216_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(KEYINPUT65), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(KEYINPUT6), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n215_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n214_), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n208_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n231_), .A2(new_n232_), .A3(G106gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n221_), .B2(new_n224_), .ZN(new_n234_));
  INV_X1    g033(.A(G85gat), .ZN(new_n235_));
  INV_X1    g034(.A(G92gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT9), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n237_), .A2(new_n238_), .B1(new_n239_), .B2(G92gat), .ZN(new_n240_));
  NOR3_X1   g039(.A1(new_n226_), .A2(new_n227_), .A3(KEYINPUT9), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT64), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n239_), .A3(new_n238_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n236_), .A2(KEYINPUT9), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n243_), .B(new_n244_), .C1(new_n228_), .C2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n234_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n212_), .A2(new_n213_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n222_), .A2(new_n223_), .A3(new_n215_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n215_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(KEYINPUT8), .A3(new_n228_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n230_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G57gat), .B(G64gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT11), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT67), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n256_), .A2(KEYINPUT11), .ZN(new_n259_));
  XOR2_X1   g058(.A(G71gat), .B(G78gat), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n258_), .B(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n230_), .A2(new_n247_), .A3(new_n252_), .A4(KEYINPUT66), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n255_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT68), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n255_), .A2(new_n262_), .A3(new_n266_), .A4(new_n263_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n255_), .A2(new_n263_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n259_), .A2(new_n260_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n258_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n265_), .A2(new_n267_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G230gat), .A2(G233gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n272_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT12), .B1(new_n268_), .B2(new_n270_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n270_), .A2(KEYINPUT12), .A3(new_n253_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n264_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n274_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n273_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n207_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n207_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n285_), .A2(new_n276_), .A3(new_n281_), .A4(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(KEYINPUT13), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT13), .B1(new_n284_), .B2(new_n287_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n202_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n289_), .A2(new_n290_), .A3(new_n202_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT77), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G15gat), .B(G22gat), .ZN(new_n297_));
  INV_X1    g096(.A(G1gat), .ZN(new_n298_));
  INV_X1    g097(.A(G8gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT14), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n295_), .A2(KEYINPUT77), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n295_), .A2(KEYINPUT77), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n303_), .A2(new_n300_), .A3(new_n297_), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT78), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n306_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(new_n270_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G127gat), .B(G155gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT16), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G183gat), .B(G211gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT17), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n315_), .A2(new_n316_), .ZN(new_n318_));
  OR3_X1    g117(.A1(new_n311_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n311_), .A2(new_n317_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT36), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G190gat), .B(G218gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G134gat), .B(G162gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G29gat), .B(G36gat), .Z(new_n326_));
  XOR2_X1   g125(.A(G43gat), .B(G50gat), .Z(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G29gat), .B(G36gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G43gat), .B(G50gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n255_), .A2(new_n332_), .A3(new_n263_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n328_), .A2(KEYINPUT15), .A3(new_n331_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT15), .B1(new_n328_), .B2(new_n331_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n253_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G232gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT34), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n339_), .A2(KEYINPUT35), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(KEYINPUT35), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n333_), .A2(new_n337_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(KEYINPUT72), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n253_), .A2(new_n336_), .A3(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n333_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n347_), .A2(KEYINPUT73), .A3(new_n340_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT73), .B1(new_n347_), .B2(new_n340_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n325_), .B(new_n343_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n351_), .B(new_n343_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n325_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n322_), .A2(new_n350_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n352_), .A2(new_n322_), .A3(new_n353_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(new_n356_), .B2(KEYINPUT37), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n350_), .A2(new_n322_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n352_), .A2(new_n353_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n352_), .A2(new_n322_), .A3(new_n353_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT37), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(KEYINPUT37), .A3(new_n361_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n360_), .A2(KEYINPUT75), .A3(KEYINPUT37), .A4(new_n361_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n357_), .A2(new_n365_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n294_), .A2(new_n321_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT23), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT24), .ZN(new_n376_));
  INV_X1    g175(.A(G169gat), .ZN(new_n377_));
  INV_X1    g176(.A(G176gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT25), .B(G183gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT26), .B(G190gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n381_), .A2(new_n382_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n380_), .A2(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n375_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(G169gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G15gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n395_), .B(KEYINPUT30), .Z(new_n396_));
  XNOR2_X1  g195(.A(new_n393_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT81), .B(G43gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G127gat), .B(G134gat), .Z(new_n400_));
  XOR2_X1   g199(.A(G113gat), .B(G120gat), .Z(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G127gat), .B(G134gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G113gat), .B(G120gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(KEYINPUT82), .A3(new_n405_), .ZN(new_n406_));
  OR3_X1    g205(.A1(new_n403_), .A2(new_n404_), .A3(KEYINPUT82), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT31), .ZN(new_n409_));
  XOR2_X1   g208(.A(G71gat), .B(G99gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n399_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n399_), .A2(new_n411_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT1), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT1), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(G155gat), .A3(G162gat), .ZN(new_n420_));
  OR2_X1    g219(.A1(G155gat), .A2(G162gat), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .A4(KEYINPUT83), .ZN(new_n422_));
  OR3_X1    g221(.A1(new_n417_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n423_));
  XOR2_X1   g222(.A(G141gat), .B(G148gat), .Z(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT3), .ZN(new_n426_));
  INV_X1    g225(.A(G141gat), .ZN(new_n427_));
  INV_X1    g226(.A(G148gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G141gat), .A2(G148gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT2), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n429_), .A2(new_n432_), .A3(new_n433_), .A4(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n421_), .A2(new_n417_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n425_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n425_), .A2(new_n437_), .A3(KEYINPUT84), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT29), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT85), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n440_), .A2(new_n445_), .A3(KEYINPUT29), .A4(new_n441_), .ZN(new_n446_));
  OR2_X1    g245(.A1(G197gat), .A2(G204gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT87), .B(G197gat), .ZN(new_n448_));
  INV_X1    g247(.A(G204gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT21), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT89), .ZN(new_n453_));
  XOR2_X1   g252(.A(G211gat), .B(G218gat), .Z(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n449_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n451_), .B1(G197gat), .B2(G204gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n454_), .B1(new_n457_), .B2(KEYINPUT88), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n455_), .A2(new_n459_), .A3(new_n456_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n450_), .A2(new_n461_), .A3(new_n451_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n453_), .A2(new_n458_), .A3(new_n460_), .A4(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT90), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n450_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n450_), .A2(new_n464_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(KEYINPUT21), .A3(new_n466_), .A4(new_n454_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(G228gat), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n444_), .A2(new_n446_), .A3(new_n468_), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(KEYINPUT91), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT91), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n463_), .A2(new_n474_), .A3(new_n467_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n473_), .A2(new_n475_), .B1(KEYINPUT29), .B2(new_n438_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n416_), .B(new_n472_), .C1(new_n476_), .C2(new_n471_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n442_), .A2(new_n443_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G22gat), .B(G50gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT28), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n480_), .B(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n472_), .B1(new_n476_), .B2(new_n471_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n415_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n477_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n486_), .A2(KEYINPUT92), .A3(new_n477_), .A4(new_n483_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G225gat), .A2(G233gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n440_), .A2(new_n441_), .A3(new_n408_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT95), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT95), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n440_), .A2(new_n408_), .A3(new_n494_), .A4(new_n441_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n438_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT4), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT4), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n492_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n491_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n496_), .A2(new_n491_), .A3(new_n498_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT98), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n497_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT98), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n491_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G1gat), .B(G29gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT97), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G57gat), .B(G85gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n510_), .A2(KEYINPUT99), .A3(KEYINPUT33), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT99), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n502_), .B1(new_n506_), .B2(new_n501_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n491_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n522_), .A2(new_n517_), .A3(new_n505_), .A4(new_n508_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT33), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n519_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G8gat), .B(G36gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G64gat), .B(G92gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G226gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT19), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n393_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT22), .B(G169gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT93), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n378_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n389_), .A2(new_n385_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n540_), .A2(new_n541_), .B1(new_n380_), .B2(new_n386_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n533_), .B1(new_n536_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n463_), .A2(new_n393_), .A3(new_n467_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT20), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n542_), .B1(new_n467_), .B2(new_n463_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n533_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n531_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n547_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n551_), .A2(KEYINPUT20), .A3(new_n533_), .A4(new_n545_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n393_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n468_), .A2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n554_), .A2(KEYINPUT20), .A3(new_n543_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n552_), .B(new_n530_), .C1(new_n555_), .C2(new_n533_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n516_), .B1(new_n499_), .B2(new_n491_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n491_), .B2(new_n520_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n523_), .A2(new_n524_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n518_), .A2(new_n525_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n531_), .A2(KEYINPUT32), .ZN(new_n563_));
  INV_X1    g362(.A(new_n544_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n564_), .B2(new_n552_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n473_), .A2(new_n475_), .A3(new_n542_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n534_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n548_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n546_), .A2(new_n547_), .A3(new_n533_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n565_), .B1(new_n571_), .B2(new_n563_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n516_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n523_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n572_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n490_), .B1(new_n562_), .B2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n574_), .A2(new_n575_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n550_), .A2(KEYINPUT27), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n530_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n579_), .A2(new_n580_), .B1(new_n557_), .B2(new_n582_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n490_), .A2(new_n578_), .A3(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n414_), .B1(new_n577_), .B2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n490_), .A2(new_n414_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n578_), .A3(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT80), .B1(new_n306_), .B2(new_n332_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n306_), .A2(new_n332_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n336_), .A2(new_n305_), .A3(new_n302_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n306_), .A2(new_n332_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595_));
  MUX2_X1   g394(.A(new_n591_), .B(new_n594_), .S(new_n595_), .Z(new_n596_));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G169gat), .B(G197gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n596_), .B(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n588_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n373_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT102), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT38), .ZN(new_n606_));
  AOI211_X1 g405(.A(G1gat), .B(new_n578_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n604_), .A2(KEYINPUT102), .A3(KEYINPUT38), .A4(new_n607_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n601_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n294_), .A2(new_n611_), .A3(new_n321_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n588_), .A2(new_n356_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(KEYINPUT103), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n588_), .B2(new_n356_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT104), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT104), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n612_), .B(new_n619_), .C1(new_n614_), .C2(new_n616_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n578_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n609_), .B(new_n610_), .C1(new_n298_), .C2(new_n621_), .ZN(G1324gat));
  XNOR2_X1  g421(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n613_), .B(KEYINPUT103), .ZN(new_n624_));
  INV_X1    g423(.A(new_n583_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n612_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n626_), .A2(new_n627_), .A3(G8gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n626_), .B2(G8gat), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n604_), .A2(new_n299_), .A3(new_n625_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n623_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n631_), .B(new_n623_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1325gat));
  INV_X1    g434(.A(new_n414_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n619_), .B1(new_n624_), .B2(new_n612_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n620_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT106), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n640_), .A3(G15gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n414_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n642_));
  INV_X1    g441(.A(G15gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT106), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n641_), .A2(new_n644_), .A3(KEYINPUT41), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n604_), .A2(new_n643_), .A3(new_n636_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT107), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n648_), .A3(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n604_), .A2(new_n652_), .A3(new_n490_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n490_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n655_), .A2(new_n652_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n656_), .A2(KEYINPUT42), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(KEYINPUT42), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n653_), .B1(new_n657_), .B2(new_n658_), .ZN(G1327gat));
  NOR2_X1   g458(.A1(new_n294_), .A2(new_n611_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n321_), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n356_), .B(new_n661_), .C1(new_n585_), .C2(new_n587_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n578_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G29gat), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n370_), .B2(KEYINPUT108), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n588_), .A2(new_n370_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n588_), .B(new_n370_), .C1(KEYINPUT108), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n293_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n291_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(new_n601_), .A3(new_n321_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT44), .B1(new_n672_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  AOI211_X1 g477(.A(new_n678_), .B(new_n675_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n665_), .A2(G29gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n666_), .B1(new_n680_), .B2(new_n681_), .ZN(G1328gat));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n664_), .A2(new_n683_), .A3(new_n625_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n684_), .B(new_n685_), .Z(new_n686_));
  NAND2_X1  g485(.A1(new_n672_), .A2(new_n676_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n678_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n676_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G36gat), .B1(new_n690_), .B2(new_n583_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n686_), .A2(new_n691_), .A3(KEYINPUT110), .A4(new_n692_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n692_), .A2(KEYINPUT110), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(KEYINPUT110), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n683_), .B1(new_n680_), .B2(new_n625_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n684_), .B(new_n685_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n694_), .B(new_n695_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n693_), .A2(new_n698_), .ZN(G1329gat));
  INV_X1    g498(.A(G43gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n700_), .B1(new_n663_), .B2(new_n414_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT111), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n636_), .A2(G43gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n690_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g504(.A(KEYINPUT113), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n688_), .A2(new_n707_), .A3(new_n490_), .A4(new_n689_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G50gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n680_), .B2(new_n490_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n688_), .A2(new_n490_), .A3(new_n689_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT112), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n713_), .A2(KEYINPUT113), .A3(G50gat), .A4(new_n708_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n654_), .A2(G50gat), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT114), .Z(new_n717_));
  NAND2_X1  g516(.A1(new_n664_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1331gat));
  INV_X1    g518(.A(G57gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n674_), .A2(new_n601_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n624_), .A2(new_n661_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(new_n665_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n370_), .A2(new_n321_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n721_), .A2(new_n588_), .A3(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n725_), .A2(new_n720_), .A3(new_n665_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1332gat));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n728_), .A3(new_n625_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n722_), .A2(new_n625_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G64gat), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT48), .B(new_n728_), .C1(new_n722_), .C2(new_n625_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(G1333gat));
  INV_X1    g533(.A(G71gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n725_), .A2(new_n735_), .A3(new_n636_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT49), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n722_), .A2(new_n636_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(G71gat), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT49), .B(new_n735_), .C1(new_n722_), .C2(new_n636_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1334gat));
  INV_X1    g540(.A(G78gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n725_), .A2(new_n742_), .A3(new_n490_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n722_), .A2(new_n490_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(G78gat), .ZN(new_n746_));
  AOI211_X1 g545(.A(KEYINPUT50), .B(new_n742_), .C1(new_n722_), .C2(new_n490_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(G1335gat));
  NAND2_X1  g547(.A1(new_n721_), .A2(new_n321_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n751_), .A2(new_n235_), .A3(new_n578_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n721_), .A2(new_n662_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n665_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n754_), .A2(KEYINPUT115), .A3(new_n235_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT115), .B1(new_n754_), .B2(new_n235_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n752_), .A2(new_n755_), .A3(new_n756_), .ZN(G1336gat));
  OAI21_X1  g556(.A(G92gat), .B1(new_n751_), .B2(new_n583_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n753_), .A2(new_n236_), .A3(new_n625_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1337gat));
  OAI21_X1  g559(.A(G99gat), .B1(new_n751_), .B2(new_n414_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n414_), .A2(new_n232_), .A3(new_n231_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n753_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g564(.A1(new_n753_), .A2(new_n211_), .A3(new_n490_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n750_), .A2(new_n490_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G106gat), .ZN(new_n769_));
  AOI211_X1 g568(.A(KEYINPUT52), .B(new_n211_), .C1(new_n750_), .C2(new_n490_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n262_), .B1(new_n255_), .B2(new_n263_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n264_), .B(new_n278_), .C1(new_n774_), .C2(KEYINPUT12), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n775_), .B2(new_n275_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT117), .B1(new_n280_), .B2(new_n274_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n775_), .A2(new_n778_), .A3(new_n275_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT55), .B1(new_n280_), .B2(new_n274_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n775_), .B2(new_n275_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n280_), .A2(KEYINPUT117), .A3(new_n274_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n780_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n207_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT118), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n207_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n785_), .A2(new_n791_), .A3(KEYINPUT56), .A4(new_n207_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n787_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n596_), .A2(new_n600_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n591_), .A2(new_n595_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n594_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n795_), .B(new_n600_), .C1(new_n595_), .C2(new_n796_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n287_), .A2(new_n794_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n793_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n793_), .A2(KEYINPUT58), .A3(new_n798_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n370_), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n601_), .A2(new_n287_), .A3(KEYINPUT116), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n601_), .A2(new_n287_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n785_), .B2(new_n207_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n789_), .B(new_n286_), .C1(new_n780_), .C2(new_n784_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n804_), .B(new_n807_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n284_), .A2(new_n287_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(new_n794_), .A3(new_n797_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n356_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n356_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n813_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n356_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n803_), .A2(new_n816_), .A3(new_n819_), .A4(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n321_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n370_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n289_), .A2(new_n290_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n611_), .A4(new_n661_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT54), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n724_), .A2(new_n827_), .A3(new_n611_), .A4(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n822_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n586_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n831_), .A2(new_n578_), .A3(new_n625_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(G113gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n601_), .B2(KEYINPUT121), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(KEYINPUT121), .B2(new_n836_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(KEYINPUT120), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n835_), .B(new_n838_), .C1(new_n833_), .C2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n836_), .B1(new_n833_), .B2(new_n611_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1340gat));
  OAI21_X1  g642(.A(new_n835_), .B1(new_n833_), .B2(new_n840_), .ZN(new_n844_));
  OAI21_X1  g643(.A(G120gat), .B1(new_n844_), .B2(new_n674_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n833_), .ZN(new_n846_));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n674_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n846_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n847_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n845_), .A2(new_n849_), .ZN(G1341gat));
  OAI21_X1  g649(.A(G127gat), .B1(new_n844_), .B2(new_n321_), .ZN(new_n851_));
  OR3_X1    g650(.A1(new_n833_), .A2(G127gat), .A3(new_n321_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1342gat));
  OAI21_X1  g652(.A(G134gat), .B1(new_n844_), .B2(new_n823_), .ZN(new_n854_));
  OR3_X1    g653(.A1(new_n833_), .A2(G134gat), .A3(new_n356_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1343gat));
  NAND4_X1  g655(.A1(new_n665_), .A2(new_n490_), .A3(new_n583_), .A4(new_n414_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT122), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n830_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n611_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n427_), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n674_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n428_), .ZN(G1345gat));
  NOR2_X1   g662(.A1(new_n859_), .A2(new_n321_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT61), .B(G155gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  OAI21_X1  g665(.A(G162gat), .B1(new_n859_), .B2(new_n823_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n356_), .A2(G162gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n859_), .B2(new_n868_), .ZN(G1347gat));
  AOI22_X1  g668(.A1(new_n821_), .A2(new_n321_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n831_), .A2(new_n665_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NOR4_X1   g671(.A1(new_n870_), .A2(new_n583_), .A3(new_n611_), .A4(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT123), .B1(new_n873_), .B2(new_n377_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n830_), .A2(new_n625_), .A3(new_n871_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n875_), .B(G169gat), .C1(new_n876_), .C2(new_n611_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n877_), .A3(KEYINPUT62), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  OAI211_X1 g678(.A(KEYINPUT123), .B(new_n879_), .C1(new_n873_), .C2(new_n377_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n873_), .A2(new_n539_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n880_), .A3(new_n881_), .ZN(G1348gat));
  INV_X1    g681(.A(new_n876_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT124), .B(G176gat), .Z(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n294_), .A3(new_n884_), .ZN(new_n885_));
  OAI22_X1  g684(.A1(new_n876_), .A2(new_n674_), .B1(KEYINPUT124), .B2(new_n378_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1349gat));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n661_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(G183gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n381_), .B1(KEYINPUT125), .B2(G183gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n888_), .B2(new_n891_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n876_), .B2(new_n823_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n362_), .A2(new_n382_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n876_), .B2(new_n894_), .ZN(G1351gat));
  NOR3_X1   g694(.A1(new_n654_), .A2(new_n665_), .A3(new_n636_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT126), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n870_), .A2(new_n583_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n601_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n294_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n661_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT63), .B(G211gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n904_), .B2(new_n907_), .ZN(G1354gat));
  NOR2_X1   g707(.A1(new_n356_), .A2(G218gat), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n830_), .A2(new_n625_), .A3(new_n897_), .A4(new_n909_), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n870_), .A2(new_n583_), .A3(new_n823_), .A4(new_n898_), .ZN(new_n911_));
  INV_X1    g710(.A(G218gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


