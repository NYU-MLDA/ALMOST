//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205_));
  INV_X1    g004(.A(G15gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n204_), .B(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G183gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT25), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT25), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G183gat), .ZN(new_n220_));
  INV_X1    g019(.A(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT26), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT26), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G190gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n218_), .A2(new_n220_), .A3(new_n222_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n213_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n225_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n216_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n234_), .B(new_n209_), .C1(G183gat), .C2(G190gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n236_));
  OR3_X1    g035(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n208_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n241_), .A2(new_n242_), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n246_), .A2(KEYINPUT83), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(KEYINPUT83), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n246_), .A2(KEYINPUT83), .ZN(new_n252_));
  INV_X1    g051(.A(G134gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G127gat), .ZN(new_n254_));
  INV_X1    g053(.A(G127gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G134gat), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n254_), .A2(new_n256_), .A3(KEYINPUT83), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n251_), .B1(new_n252_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n250_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT31), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n245_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n245_), .A2(new_n260_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G1gat), .B(G29gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G85gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT0), .B(G57gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G141gat), .ZN(new_n269_));
  INV_X1    g068(.A(G148gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n271_), .B(new_n272_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n276_), .A2(new_n277_), .A3(KEYINPUT1), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT84), .B1(new_n275_), .B2(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n271_), .A2(new_n272_), .ZN(new_n280_));
  OR2_X1    g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT84), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(KEYINPUT1), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n280_), .A2(new_n282_), .A3(new_n283_), .A4(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n272_), .B(KEYINPUT2), .ZN(new_n287_));
  OAI22_X1  g086(.A1(KEYINPUT85), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n271_), .A2(KEYINPUT85), .A3(KEYINPUT3), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n276_), .A2(new_n277_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n286_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n259_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n286_), .A2(new_n294_), .A3(new_n250_), .A4(new_n258_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(KEYINPUT4), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G225gat), .A2(G233gat), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n286_), .A2(new_n294_), .B1(new_n250_), .B2(new_n258_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n302_), .A3(KEYINPUT97), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n296_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT97), .B1(new_n298_), .B2(new_n302_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n268_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n306_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n308_), .A2(new_n267_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n295_), .A2(KEYINPUT29), .ZN(new_n311_));
  INV_X1    g110(.A(G204gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G197gat), .ZN(new_n313_));
  INV_X1    g112(.A(G197gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G204gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT86), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(new_n314_), .B2(G204gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(KEYINPUT21), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT21), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n313_), .B(new_n315_), .C1(new_n317_), .C2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G218gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G211gat), .ZN(new_n323_));
  INV_X1    g122(.A(G211gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G218gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n319_), .A2(new_n321_), .A3(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n316_), .A2(new_n326_), .A3(KEYINPUT21), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT87), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n320_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(new_n326_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n330_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT88), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT88), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n328_), .A2(new_n330_), .A3(new_n336_), .A4(new_n333_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G228gat), .A2(G233gat), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n311_), .A2(new_n335_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n286_), .B2(new_n294_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n334_), .ZN(new_n342_));
  OAI211_X1 g141(.A(G228gat), .B(G233gat), .C1(new_n341_), .C2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G78gat), .B(G106gat), .Z(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT28), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n279_), .A2(new_n285_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(new_n340_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n347_), .A3(new_n340_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G22gat), .B(G50gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n351_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n352_), .B1(new_n355_), .B2(new_n349_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n345_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n339_), .A2(new_n343_), .A3(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n346_), .A2(new_n354_), .A3(new_n356_), .A4(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n354_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n339_), .A2(new_n357_), .A3(new_n343_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n357_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n335_), .A2(new_n337_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n238_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n225_), .A2(new_n228_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT80), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n225_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n372_), .B1(new_n376_), .B2(new_n216_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n370_), .B1(new_n371_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n227_), .B(KEYINPUT94), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT22), .B(G169gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT95), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n235_), .B(new_n379_), .C1(new_n382_), .C2(G176gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT90), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n219_), .A2(G183gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n217_), .A2(KEYINPUT25), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n222_), .A2(new_n224_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n218_), .A2(new_n220_), .A3(KEYINPUT90), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT91), .B1(new_n227_), .B2(KEYINPUT24), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(new_n213_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n227_), .A2(KEYINPUT91), .A3(KEYINPUT24), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n394_), .A3(KEYINPUT92), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT93), .B1(new_n212_), .B2(new_n215_), .ZN(new_n396_));
  AND4_X1   g195(.A1(KEYINPUT93), .A2(new_n234_), .A3(new_n215_), .A4(new_n209_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT92), .B1(new_n390_), .B2(new_n394_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n383_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n334_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n369_), .B1(new_n378_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n239_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n342_), .B(new_n383_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(KEYINPUT20), .A4(new_n369_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G64gat), .B(G92gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n403_), .A2(new_n407_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  AND4_X1   g213(.A1(new_n332_), .A2(new_n316_), .A3(new_n326_), .A4(KEYINPUT21), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n332_), .B1(new_n331_), .B2(new_n326_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n336_), .B1(new_n417_), .B2(new_n328_), .ZN(new_n418_));
  AND4_X1   g217(.A1(new_n336_), .A2(new_n328_), .A3(new_n330_), .A4(new_n333_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n377_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT20), .ZN(new_n421_));
  INV_X1    g220(.A(new_n400_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n395_), .A3(new_n398_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n342_), .B1(new_n423_), .B2(new_n383_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n368_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n414_), .B1(new_n425_), .B2(new_n406_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n365_), .B1(new_n413_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n404_), .A2(new_n405_), .A3(KEYINPUT20), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n368_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n402_), .A2(KEYINPUT20), .A3(new_n420_), .A4(new_n369_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n412_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n425_), .A2(new_n414_), .A3(new_n406_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT27), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  NOR4_X1   g234(.A1(new_n263_), .A2(new_n310_), .A3(new_n364_), .A4(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n307_), .A2(new_n309_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n427_), .A2(new_n437_), .A3(new_n364_), .A4(new_n434_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT102), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n359_), .A2(new_n363_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(new_n310_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n442_), .A2(KEYINPUT102), .A3(new_n427_), .A4(new_n434_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n305_), .A2(new_n268_), .A3(new_n306_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n296_), .A2(G225gat), .A3(G233gat), .A4(new_n297_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n446_), .A2(new_n268_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n298_), .B(new_n299_), .C1(KEYINPUT4), .C2(new_n296_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT99), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT99), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n445_), .A2(KEYINPUT33), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n309_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT98), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n412_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n433_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT98), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n309_), .A2(new_n460_), .A3(new_n454_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n453_), .A2(new_n456_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n414_), .A2(KEYINPUT32), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n307_), .A2(new_n309_), .B1(new_n464_), .B2(new_n431_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n403_), .A2(new_n407_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(KEYINPUT100), .A3(new_n463_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT100), .B1(new_n466_), .B2(new_n463_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n465_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n364_), .B1(new_n462_), .B2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n263_), .B1(new_n444_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT103), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT103), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n474_), .B(new_n263_), .C1(new_n444_), .C2(new_n471_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n436_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G57gat), .B(G64gat), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n479_));
  XOR2_X1   g278(.A(G71gat), .B(G78gat), .Z(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n479_), .A2(new_n480_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484_));
  INV_X1    g283(.A(G1gat), .ZN(new_n485_));
  INV_X1    g284(.A(G8gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G1gat), .B(G8gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n483_), .B(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G231gat), .A2(G233gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  XOR2_X1   g292(.A(G127gat), .B(G155gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(G183gat), .B(G211gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT17), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n493_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n493_), .A2(KEYINPUT17), .A3(new_n498_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G85gat), .ZN(new_n503_));
  INV_X1    g302(.A(G92gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT9), .ZN(new_n506_));
  NOR2_X1   g305(.A1(G85gat), .A2(G92gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n506_), .B1(new_n507_), .B2(KEYINPUT64), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n505_), .A2(KEYINPUT9), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n508_), .B(new_n509_), .C1(KEYINPUT64), .C2(new_n506_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT10), .B(G99gat), .Z(new_n514_));
  INV_X1    g313(.A(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n510_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT67), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n521_), .A2(G99gat), .A3(G106gat), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT7), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n513_), .B(new_n525_), .C1(new_n524_), .C2(new_n522_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n505_), .A2(new_n507_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT8), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT8), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n518_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G29gat), .B(G36gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT71), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G43gat), .B(G50gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT35), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT34), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n532_), .A2(new_n536_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT15), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n536_), .B(new_n542_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n543_), .A2(new_n532_), .A3(KEYINPUT72), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n545_));
  INV_X1    g344(.A(new_n531_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n530_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n517_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n536_), .B(KEYINPUT15), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n545_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n541_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n540_), .A2(new_n537_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT72), .B1(new_n543_), .B2(new_n532_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n548_), .A2(new_n549_), .A3(new_n545_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n552_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n541_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G190gat), .B(G218gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT74), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n553_), .A2(new_n558_), .A3(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n561_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n565_), .B1(new_n569_), .B2(KEYINPUT76), .ZN(new_n570_));
  INV_X1    g369(.A(new_n558_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n557_), .B1(new_n556_), .B2(new_n541_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n567_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT76), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT37), .B1(new_n570_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(new_n577_), .A3(new_n565_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n578_), .A2(KEYINPUT77), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT77), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n581_), .B(KEYINPUT37), .C1(new_n570_), .C2(new_n575_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n476_), .A2(new_n502_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n483_), .B(new_n517_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT12), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n532_), .A2(new_n483_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n532_), .A2(KEYINPUT12), .A3(new_n483_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n585_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n483_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n548_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT68), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n586_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n585_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n532_), .A2(KEYINPUT68), .A3(new_n483_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n591_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT5), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n599_), .A2(new_n603_), .ZN(new_n606_));
  OAI22_X1  g405(.A1(new_n605_), .A2(new_n606_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n604_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT70), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(KEYINPUT70), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n536_), .B(new_n490_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G229gat), .A2(G233gat), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n536_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(new_n490_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n549_), .B2(new_n490_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n618_), .B1(new_n621_), .B2(new_n617_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G169gat), .B(G197gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  NOR2_X1   g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(new_n625_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT79), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT79), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n622_), .A2(new_n629_), .A3(new_n625_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n626_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n615_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n584_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n437_), .B(KEYINPUT104), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n633_), .A2(G1gat), .A3(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n635_), .A2(KEYINPUT38), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(KEYINPUT38), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n573_), .A2(new_n565_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n502_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n473_), .A2(new_n475_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n436_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n631_), .ZN(new_n644_));
  AND4_X1   g443(.A1(new_n640_), .A2(new_n643_), .A3(new_n644_), .A4(new_n612_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(new_n310_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n636_), .B(new_n637_), .C1(new_n485_), .C2(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n435_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n649_), .B2(G8gat), .ZN(new_n650_));
  AOI211_X1 g449(.A(KEYINPUT39), .B(new_n486_), .C1(new_n645_), .C2(new_n435_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n435_), .A2(new_n486_), .ZN(new_n652_));
  OAI22_X1  g451(.A1(new_n650_), .A2(new_n651_), .B1(new_n633_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n653_), .B(new_n654_), .Z(G1325gat));
  INV_X1    g454(.A(new_n263_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n206_), .B1(new_n645_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT41), .ZN(new_n658_));
  INV_X1    g457(.A(new_n633_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n206_), .A3(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(G1326gat));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n645_), .B2(new_n364_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT42), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n659_), .A2(new_n662_), .A3(new_n364_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n502_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n638_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n643_), .A2(new_n644_), .A3(new_n612_), .A4(new_n668_), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n669_), .A2(KEYINPUT109), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(KEYINPUT109), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(G29gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n310_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n580_), .A2(new_n582_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n476_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n675_), .B(KEYINPUT43), .C1(new_n476_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n612_), .A2(new_n502_), .A3(new_n644_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT106), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n634_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n684_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n690_), .A2(KEYINPUT108), .A3(G29gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT108), .B1(new_n690_), .B2(G29gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n674_), .B1(new_n691_), .B2(new_n692_), .ZN(G1328gat));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(KEYINPUT46), .ZN(new_n695_));
  INV_X1    g494(.A(G36gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT44), .B1(new_n681_), .B2(new_n684_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n686_), .B(new_n683_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n696_), .B1(new_n699_), .B2(new_n435_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n435_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(G36gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n670_), .A2(new_n671_), .A3(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n704_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n670_), .A2(new_n671_), .A3(new_n706_), .A4(new_n702_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n695_), .B1(new_n700_), .B2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n687_), .A2(new_n435_), .A3(new_n689_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n705_), .A2(new_n707_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n695_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n709_), .A2(new_n714_), .ZN(G1329gat));
  NAND4_X1  g514(.A1(new_n687_), .A2(G43gat), .A3(new_n656_), .A4(new_n689_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n670_), .A2(new_n656_), .A3(new_n671_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n203_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT47), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n716_), .A2(new_n721_), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n672_), .B2(new_n364_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n364_), .A2(G50gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n699_), .B2(new_n725_), .ZN(G1331gat));
  NOR2_X1   g525(.A1(new_n612_), .A2(new_n644_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n584_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G57gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n688_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n615_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n731_), .A2(new_n476_), .A3(new_n644_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n732_), .A2(new_n310_), .A3(new_n640_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n730_), .B1(new_n733_), .B2(new_n729_), .ZN(G1332gat));
  INV_X1    g533(.A(G64gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n728_), .A2(new_n735_), .A3(new_n435_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(new_n640_), .A3(new_n435_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(G64gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G64gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1333gat));
  INV_X1    g540(.A(G71gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n728_), .A2(new_n742_), .A3(new_n656_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n732_), .A2(new_n640_), .A3(new_n656_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(new_n745_), .A3(G71gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(G71gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(G1334gat));
  INV_X1    g547(.A(G78gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n728_), .A2(new_n749_), .A3(new_n364_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n732_), .A2(new_n640_), .A3(new_n364_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(G78gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n751_), .B2(G78gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(G1335gat));
  NAND2_X1  g554(.A1(new_n727_), .A2(new_n502_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n503_), .B1(new_n757_), .B2(new_n310_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n732_), .A2(new_n668_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n759_), .A2(G85gat), .A3(new_n634_), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1336gat));
  OAI21_X1  g560(.A(new_n504_), .B1(new_n759_), .B2(new_n701_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT112), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n701_), .A2(new_n504_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n757_), .B2(new_n764_), .ZN(G1337gat));
  INV_X1    g564(.A(new_n756_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n681_), .A2(new_n656_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(G99gat), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n767_), .B2(G99gat), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT114), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n656_), .A2(new_n514_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n759_), .A2(new_n775_), .B1(KEYINPUT114), .B2(new_n772_), .ZN(new_n776_));
  NOR4_X1   g575(.A1(new_n770_), .A2(new_n771_), .A3(new_n774_), .A4(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n767_), .A2(G99gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n778_), .B2(KEYINPUT113), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n773_), .B1(new_n779_), .B2(new_n769_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1338gat));
  AOI211_X1 g580(.A(KEYINPUT52), .B(new_n515_), .C1(new_n757_), .C2(new_n364_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n681_), .A2(new_n364_), .A3(new_n766_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(G106gat), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n364_), .A2(new_n515_), .ZN(new_n786_));
  OAI22_X1  g585(.A1(new_n782_), .A2(new_n785_), .B1(new_n759_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789_));
  OAI221_X1 g588(.A(new_n789_), .B1(new_n759_), .B2(new_n786_), .C1(new_n782_), .C2(new_n785_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1339gat));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n631_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n607_), .B2(new_n611_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n580_), .A2(new_n795_), .A3(new_n667_), .A4(new_n582_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800_));
  INV_X1    g599(.A(new_n590_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n593_), .A2(KEYINPUT12), .A3(new_n586_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n596_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n800_), .B1(new_n803_), .B2(KEYINPUT55), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n591_), .A2(KEYINPUT116), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(KEYINPUT55), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n801_), .A2(new_n802_), .A3(new_n596_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n804_), .A2(new_n806_), .A3(new_n807_), .A4(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n603_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n644_), .A2(new_n608_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT117), .B1(new_n809_), .B2(new_n603_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n608_), .A2(new_n604_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n628_), .A2(new_n630_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n617_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n621_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n625_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n821_), .B(new_n822_), .C1(new_n820_), .C2(new_n616_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n819_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT118), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n819_), .A2(new_n826_), .A3(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n814_), .A2(new_n817_), .B1(new_n818_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n799_), .B1(new_n829_), .B2(new_n639_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n818_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n810_), .A2(new_n811_), .A3(KEYINPUT56), .ZN(new_n832_));
  INV_X1    g631(.A(new_n815_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n816_), .A2(KEYINPUT56), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(KEYINPUT57), .A3(new_n638_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n606_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n810_), .A2(KEYINPUT56), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n809_), .A2(new_n813_), .A3(new_n603_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n838_), .A2(new_n839_), .A3(KEYINPUT58), .A4(new_n840_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n583_), .A3(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n830_), .A2(new_n837_), .A3(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n798_), .B1(new_n846_), .B2(new_n502_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n688_), .A2(new_n701_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n848_), .A2(new_n263_), .A3(new_n364_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n644_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT120), .B1(new_n853_), .B2(KEYINPUT119), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n836_), .A2(new_n638_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n841_), .A2(new_n842_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n855_), .A2(new_n799_), .B1(new_n856_), .B2(new_n844_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n667_), .B1(new_n857_), .B2(new_n837_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n849_), .B(new_n854_), .C1(new_n858_), .C2(new_n798_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n849_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n853_), .B1(new_n847_), .B2(new_n862_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n859_), .A2(new_n863_), .A3(KEYINPUT121), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT121), .B1(new_n859_), .B2(new_n863_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n644_), .A2(G113gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n852_), .B1(new_n866_), .B2(new_n867_), .ZN(G1340gat));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n612_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n851_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n869_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n731_), .B1(new_n859_), .B2(new_n863_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n869_), .ZN(G1341gat));
  AOI21_X1  g672(.A(G127gat), .B1(new_n851_), .B2(new_n667_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n502_), .A2(new_n255_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n866_), .B2(new_n875_), .ZN(G1342gat));
  INV_X1    g675(.A(new_n847_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n639_), .A3(new_n849_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(KEYINPUT122), .A3(new_n253_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n847_), .A2(new_n638_), .A3(new_n850_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(G134gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n676_), .A2(new_n253_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n866_), .B2(new_n884_), .ZN(G1343gat));
  NOR2_X1   g684(.A1(new_n847_), .A2(new_n656_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n848_), .A2(new_n441_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n631_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n269_), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n731_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n270_), .ZN(G1345gat));
  NOR2_X1   g691(.A1(new_n888_), .A2(new_n502_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT61), .B(G155gat), .Z(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n888_), .B2(new_n676_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n638_), .A2(G162gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n888_), .B2(new_n897_), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n263_), .A2(new_n364_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n435_), .A3(new_n634_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n847_), .A2(new_n631_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(G169gat), .ZN(new_n904_));
  INV_X1    g703(.A(G169gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT123), .B1(new_n901_), .B2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n904_), .A2(KEYINPUT62), .A3(new_n906_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n902_), .A2(new_n382_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT123), .B(new_n909_), .C1(new_n901_), .C2(new_n905_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n907_), .A2(new_n908_), .A3(new_n910_), .ZN(G1348gat));
  NOR2_X1   g710(.A1(new_n847_), .A2(new_n900_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  OR3_X1    g712(.A1(new_n913_), .A2(G176gat), .A3(new_n612_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G176gat), .B1(new_n913_), .B2(new_n731_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1349gat));
  NAND2_X1  g715(.A1(new_n912_), .A2(new_n667_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n217_), .B2(new_n917_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n913_), .B2(new_n676_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n912_), .A2(new_n639_), .A3(new_n388_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1351gat));
  AND2_X1   g721(.A1(new_n435_), .A2(new_n442_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n886_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n631_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n314_), .ZN(G1352gat));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n731_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT124), .B(G204gat), .Z(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1353gat));
  INV_X1    g728(.A(new_n924_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n931_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n932_));
  AOI211_X1 g731(.A(new_n932_), .B(new_n502_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n930_), .A2(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n931_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n930_), .A2(new_n933_), .A3(new_n935_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1354gat));
  AND3_X1   g738(.A1(new_n886_), .A2(new_n639_), .A3(new_n923_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  AOI21_X1  g740(.A(G218gat), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(KEYINPUT126), .B1(new_n924_), .B2(new_n638_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n583_), .A2(G218gat), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(KEYINPUT127), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n942_), .A2(new_n943_), .B1(new_n930_), .B2(new_n945_), .ZN(G1355gat));
endmodule


