//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_;
  XNOR2_X1  g000(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT24), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(new_n214_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT25), .B(G183gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n212_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n206_), .B2(KEYINPUT22), .ZN(new_n224_));
  AOI21_X1  g023(.A(G176gat), .B1(new_n206_), .B2(KEYINPUT22), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT22), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(KEYINPUT84), .A3(G169gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT85), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G183gat), .ZN(new_n231_));
  INV_X1    g030(.A(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n213_), .A2(new_n215_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n233_), .B(new_n234_), .C1(new_n217_), .C2(new_n213_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT85), .A4(new_n227_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n230_), .A2(new_n235_), .A3(new_n210_), .A4(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT86), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n222_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n222_), .B2(new_n237_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G197gat), .B(G204gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT90), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G211gat), .B(G218gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT21), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT21), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n244_), .A2(new_n248_), .A3(new_n245_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT91), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n242_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n245_), .B1(new_n250_), .B2(new_n242_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n247_), .A2(new_n249_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n240_), .A2(new_n241_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n234_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n217_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(new_n214_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n212_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT93), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n220_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n220_), .A2(new_n259_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n219_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n218_), .A2(new_n233_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n210_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT22), .B(G169gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n264_), .B1(new_n265_), .B2(new_n207_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n258_), .A2(new_n262_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n252_), .A2(new_n251_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n249_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n248_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT20), .B1(new_n267_), .B2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n205_), .B1(new_n254_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n204_), .A2(KEYINPUT20), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n262_), .A2(new_n257_), .A3(new_n212_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n263_), .A2(new_n266_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n271_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT94), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n279_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n253_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n267_), .A2(KEYINPUT94), .A3(new_n271_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n273_), .A2(new_n278_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT103), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n273_), .A2(new_n287_), .A3(KEYINPUT103), .A4(new_n278_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT27), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT20), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n280_), .A2(new_n281_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(new_n253_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n222_), .A2(new_n237_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT86), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n239_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n296_), .B(new_n204_), .C1(new_n299_), .C2(new_n253_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n285_), .A2(KEYINPUT20), .A3(new_n282_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n300_), .B1(new_n301_), .B2(new_n204_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n278_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n293_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n292_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT104), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n292_), .A2(new_n304_), .A3(KEYINPUT104), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n288_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n278_), .B1(new_n273_), .B2(new_n287_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n293_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT88), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT3), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT2), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(KEYINPUT1), .B2(new_n319_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(KEYINPUT1), .B2(new_n319_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n314_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n326_), .A2(new_n316_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n313_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n318_), .A2(new_n322_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT88), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(KEYINPUT29), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G228gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT89), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n253_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n253_), .B1(new_n338_), .B2(new_n330_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G228gat), .A3(G233gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  AOI211_X1 g140(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n329_), .C2(new_n331_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n329_), .A2(new_n331_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n338_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT28), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n341_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n344_), .B2(new_n338_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n340_), .B(new_n337_), .C1(new_n349_), .C2(new_n342_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G22gat), .B(G50gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n347_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n309_), .A2(new_n312_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G227gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(G71gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G99gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n299_), .B(new_n362_), .Z(new_n363_));
  XOR2_X1   g162(.A(G127gat), .B(G134gat), .Z(new_n364_));
  XOR2_X1   g163(.A(G113gat), .B(G120gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n363_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT87), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT30), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT31), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n368_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n363_), .B(new_n366_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n372_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n329_), .A2(new_n331_), .A3(new_n367_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n367_), .A2(KEYINPUT96), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT96), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n366_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n330_), .A3(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n379_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT100), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT100), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n379_), .A2(new_n384_), .A3(new_n387_), .A4(new_n380_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT99), .ZN(new_n391_));
  XOR2_X1   g190(.A(G1gat), .B(G29gat), .Z(new_n392_));
  OR2_X1    g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G57gat), .B(G85gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n392_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n379_), .A2(KEYINPUT4), .A3(new_n384_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n380_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT97), .B(KEYINPUT4), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n329_), .A2(new_n331_), .A3(new_n367_), .A4(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n389_), .A2(new_n399_), .A3(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n398_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n378_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n357_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n356_), .A2(new_n408_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n292_), .A2(new_n304_), .A3(KEYINPUT104), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT104), .B1(new_n292_), .B2(new_n304_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n412_), .B(new_n312_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT105), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT105), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n309_), .A2(new_n417_), .A3(new_n312_), .A4(new_n412_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT102), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n400_), .A2(new_n380_), .A3(new_n403_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n379_), .A2(new_n401_), .A3(new_n384_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(new_n398_), .A3(KEYINPUT101), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT101), .B1(new_n421_), .B2(new_n398_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n419_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n426_), .A2(KEYINPUT102), .A3(new_n420_), .A4(new_n422_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n405_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n310_), .A2(new_n311_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n389_), .A2(KEYINPUT33), .A3(new_n399_), .A4(new_n404_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n278_), .A2(KEYINPUT32), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n302_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n273_), .A2(new_n287_), .A3(new_n434_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n408_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n356_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n416_), .A2(new_n418_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n411_), .B1(new_n441_), .B2(new_n377_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G43gat), .B(G50gat), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G29gat), .B(G36gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT75), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n445_), .A2(KEYINPUT75), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n444_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(new_n446_), .A3(new_n443_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT14), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT79), .B(G1gat), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(G8gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(G15gat), .B(G22gat), .Z(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT80), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(KEYINPUT79), .A2(G1gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(KEYINPUT79), .A2(G1gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(G8gat), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT14), .ZN(new_n461_));
  INV_X1    g260(.A(new_n456_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT80), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G8gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n457_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n457_), .B2(new_n464_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n452_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G229gat), .A2(G233gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT76), .B(KEYINPUT15), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n452_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n449_), .A2(new_n451_), .A3(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n465_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n455_), .A2(KEYINPUT80), .A3(new_n456_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n463_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n466_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n469_), .B(new_n470_), .C1(new_n476_), .C2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n480_), .A2(new_n466_), .A3(new_n451_), .A4(new_n449_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n469_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n470_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT81), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT81), .ZN(new_n487_));
  AOI211_X1 g286(.A(new_n487_), .B(new_n470_), .C1(new_n469_), .C2(new_n483_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n482_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G113gat), .B(G141gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT82), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G169gat), .B(G197gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n482_), .B(new_n493_), .C1(new_n486_), .C2(new_n488_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n442_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT73), .ZN(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT6), .B1(new_n361_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(G99gat), .A3(G106gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(G85gat), .ZN(new_n506_));
  INV_X1    g305(.A(G92gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(KEYINPUT9), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT9), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(G85gat), .A3(G92gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n505_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT64), .ZN(new_n514_));
  XOR2_X1   g313(.A(KEYINPUT10), .B(G99gat), .Z(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(new_n501_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n514_), .A3(new_n501_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n513_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n520_));
  NAND2_X1  g319(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(new_n361_), .A3(new_n501_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n520_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT65), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n530_));
  NOR2_X1   g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n530_), .A2(KEYINPUT67), .A3(new_n521_), .A4(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n524_), .A2(new_n529_), .A3(new_n505_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n508_), .A2(new_n509_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT68), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT8), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT8), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n538_), .A3(new_n535_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n519_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n541_));
  XOR2_X1   g340(.A(G57gat), .B(G64gat), .Z(new_n542_));
  INV_X1    g341(.A(KEYINPUT11), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT69), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n543_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G71gat), .B(G78gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(G57gat), .B(G64gat), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(KEYINPUT11), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .A4(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n546_), .B1(KEYINPUT11), .B2(new_n547_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n547_), .A2(new_n548_), .A3(KEYINPUT11), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n547_), .B2(KEYINPUT11), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  NOR3_X1   g354(.A1(new_n540_), .A2(new_n541_), .A3(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n505_), .A2(new_n512_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n518_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n510_), .B(new_n557_), .C1(new_n558_), .C2(new_n516_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n533_), .A2(new_n538_), .A3(new_n535_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n538_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n555_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT12), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n555_), .B(new_n559_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n556_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n566_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n537_), .A2(new_n539_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n555_), .B1(new_n570_), .B2(new_n559_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n565_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n569_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT70), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n562_), .A2(new_n563_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n565_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT70), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n569_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n568_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G120gat), .B(G148gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT72), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n500_), .B1(new_n579_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n541_), .B1(new_n540_), .B2(new_n555_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n569_), .B1(new_n540_), .B2(new_n555_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n562_), .A2(KEYINPUT12), .A3(new_n563_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n577_), .B1(new_n576_), .B2(new_n569_), .ZN(new_n592_));
  AOI211_X1 g391(.A(KEYINPUT70), .B(new_n566_), .C1(new_n575_), .C2(new_n565_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n591_), .B(new_n584_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(KEYINPUT73), .A3(new_n585_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n587_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n587_), .A2(KEYINPUT13), .A3(new_n594_), .A4(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT74), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n480_), .A2(new_n466_), .A3(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n480_), .B2(new_n466_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n563_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n563_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n607_));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT17), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n606_), .A2(new_n607_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT17), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n452_), .B(new_n559_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT77), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT77), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n570_), .A2(new_n620_), .A3(new_n452_), .A4(new_n559_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT35), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT34), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI22_X1  g425(.A1(new_n475_), .A2(new_n562_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n626_), .A2(new_n623_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT78), .ZN(new_n631_));
  INV_X1    g430(.A(new_n629_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n622_), .A2(new_n632_), .A3(new_n627_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n634_), .A2(KEYINPUT36), .A3(new_n638_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n622_), .A2(new_n632_), .A3(new_n627_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n632_), .B1(new_n622_), .B2(new_n627_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n637_), .B1(new_n642_), .B2(new_n631_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n630_), .A2(new_n637_), .A3(new_n633_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT36), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n639_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT37), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n640_), .A2(new_n641_), .A3(KEYINPUT78), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n645_), .B(new_n644_), .C1(new_n649_), .C2(new_n637_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n639_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n648_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n499_), .A2(new_n602_), .A3(new_n617_), .A4(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(new_n409_), .A3(new_n454_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n655_), .A2(KEYINPUT38), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(KEYINPUT38), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n647_), .A2(KEYINPUT106), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT106), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n659_), .B(new_n639_), .C1(new_n643_), .C2(new_n646_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n442_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n617_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n601_), .A2(new_n498_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G1gat), .B1(new_n665_), .B2(new_n409_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n656_), .A2(new_n657_), .A3(new_n666_), .ZN(G1324gat));
  NAND2_X1  g466(.A1(new_n309_), .A2(new_n312_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n662_), .A2(new_n668_), .A3(new_n664_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(G8gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n669_), .B2(G8gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n668_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(G8gat), .ZN(new_n675_));
  OAI22_X1  g474(.A1(new_n672_), .A2(new_n673_), .B1(new_n654_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n676_), .B(new_n677_), .Z(G1325gat));
  NAND3_X1  g477(.A1(new_n662_), .A2(new_n378_), .A3(new_n664_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT41), .B1(new_n679_), .B2(G15gat), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n377_), .A2(G15gat), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n681_), .A2(new_n682_), .B1(new_n654_), .B2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT108), .Z(G1326gat));
  OAI21_X1  g484(.A(G22gat), .B1(new_n665_), .B2(new_n356_), .ZN(new_n686_));
  XOR2_X1   g485(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n356_), .A2(G22gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n654_), .B2(new_n689_), .ZN(G1327gat));
  NAND2_X1  g489(.A1(new_n661_), .A2(new_n663_), .ZN(new_n691_));
  NOR4_X1   g490(.A1(new_n442_), .A2(new_n498_), .A3(new_n601_), .A4(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G29gat), .B1(new_n692_), .B2(new_n408_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n442_), .B2(new_n653_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n648_), .A2(new_n652_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n415_), .A2(KEYINPUT105), .B1(new_n439_), .B2(new_n356_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n378_), .B1(new_n697_), .B2(new_n418_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n695_), .B(new_n696_), .C1(new_n698_), .C2(new_n411_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n694_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n601_), .A2(new_n498_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n663_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT44), .B1(new_n700_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n705_), .B(new_n702_), .C1(new_n694_), .C2(new_n699_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n408_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n693_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  NOR2_X1   g508(.A1(new_n674_), .A2(G36gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n692_), .A2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT45), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n704_), .A2(new_n706_), .A3(new_n674_), .ZN(new_n713_));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(KEYINPUT46), .B(new_n712_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1329gat));
  AOI21_X1  g518(.A(G43gat), .B1(new_n692_), .B2(new_n378_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n378_), .A2(G43gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n707_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(G1330gat));
  NOR2_X1   g523(.A1(new_n356_), .A2(G50gat), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT110), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n692_), .A2(new_n726_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n704_), .A2(new_n706_), .A3(new_n356_), .ZN(new_n728_));
  INV_X1    g527(.A(G50gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(G1331gat));
  NOR2_X1   g529(.A1(new_n442_), .A2(new_n497_), .ZN(new_n731_));
  AND4_X1   g530(.A1(new_n601_), .A2(new_n731_), .A3(new_n617_), .A4(new_n653_), .ZN(new_n732_));
  INV_X1    g531(.A(G57gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n408_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n602_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n617_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n662_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n739_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(new_n408_), .A3(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n734_), .B1(new_n742_), .B2(new_n733_), .ZN(G1332gat));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n732_), .A2(new_n744_), .A3(new_n668_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n668_), .A3(new_n741_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n747_), .A3(G64gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(G64gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1333gat));
  NAND3_X1  g549(.A1(new_n732_), .A2(new_n359_), .A3(new_n378_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n740_), .A2(new_n378_), .A3(new_n741_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G71gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G71gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(G1334gat));
  INV_X1    g555(.A(G78gat), .ZN(new_n757_));
  INV_X1    g556(.A(new_n356_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n732_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n740_), .A2(new_n758_), .A3(new_n741_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G78gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G78gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1335gat));
  NOR2_X1   g563(.A1(new_n602_), .A2(new_n691_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n731_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n506_), .A3(new_n408_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n601_), .A2(new_n498_), .A3(new_n663_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n694_), .B2(new_n699_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n408_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n771_), .B2(new_n506_), .ZN(G1336gat));
  NAND3_X1  g571(.A1(new_n770_), .A2(G92gat), .A3(new_n668_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n767_), .A2(new_n668_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT112), .A3(new_n507_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT112), .B1(new_n774_), .B2(new_n507_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT113), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n773_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1337gat));
  AOI21_X1  g581(.A(new_n361_), .B1(new_n770_), .B2(new_n378_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n515_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n766_), .A2(new_n377_), .A3(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g586(.A1(new_n767_), .A2(new_n501_), .A3(new_n758_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n770_), .A2(new_n758_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G106gat), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT52), .B(new_n501_), .C1(new_n770_), .C2(new_n758_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(new_n788_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  OR2_X1    g596(.A1(new_n736_), .A2(KEYINPUT114), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n736_), .A2(KEYINPUT114), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n599_), .A2(new_n798_), .A3(new_n600_), .A4(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT54), .B1(new_n696_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n601_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n798_), .A2(new_n799_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n653_), .A4(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n801_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n591_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n588_), .A2(new_n590_), .A3(new_n565_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n569_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT55), .A4(new_n590_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n585_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n495_), .A2(new_n496_), .B1(new_n579_), .B2(new_n584_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n493_), .B1(new_n484_), .B2(new_n470_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n469_), .B(new_n485_), .C1(new_n476_), .C2(new_n481_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n496_), .A2(new_n822_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n818_), .A2(new_n819_), .B1(new_n597_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n807_), .B1(new_n661_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT115), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n827_), .B(new_n807_), .C1(new_n661_), .C2(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n596_), .A2(new_n594_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT73), .B1(new_n595_), .B2(new_n585_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n823_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n585_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n819_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(KEYINPUT57), .A3(new_n660_), .A4(new_n658_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n594_), .A2(new_n496_), .A3(new_n822_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT58), .B(new_n837_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n840_), .A2(new_n652_), .A3(new_n648_), .A4(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n826_), .A2(new_n828_), .A3(new_n836_), .A4(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n806_), .B1(new_n843_), .B2(new_n663_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n357_), .A2(new_n409_), .A3(new_n377_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(G113gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n497_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n836_), .A2(new_n842_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n660_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n659_), .B1(new_n650_), .B2(new_n639_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT57), .B1(new_n853_), .B2(new_n835_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n663_), .B1(new_n850_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT116), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n801_), .A2(new_n805_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n858_), .B(new_n663_), .C1(new_n850_), .C2(new_n854_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n856_), .A2(new_n857_), .A3(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n846_), .A2(KEYINPUT59), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT117), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(new_n864_), .A3(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT59), .B1(new_n844_), .B2(new_n846_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n497_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n849_), .B1(new_n869_), .B2(new_n848_), .ZN(G1340gat));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n867_), .A2(new_n735_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n866_), .B2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n802_), .A2(KEYINPUT60), .ZN(new_n874_));
  MUX2_X1   g673(.A(KEYINPUT60), .B(new_n874_), .S(new_n871_), .Z(new_n875_));
  NAND2_X1  g674(.A1(new_n847_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT118), .B1(new_n873_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n867_), .A2(new_n735_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n879_), .B(new_n876_), .C1(new_n881_), .C2(new_n871_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n882_), .ZN(G1341gat));
  INV_X1    g682(.A(G127gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n847_), .A2(new_n884_), .A3(new_n617_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n866_), .A2(new_n617_), .A3(new_n867_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n887_), .B2(new_n884_), .ZN(G1342gat));
  XOR2_X1   g687(.A(KEYINPUT119), .B(G134gat), .Z(new_n889_));
  NOR2_X1   g688(.A1(new_n653_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n865_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n864_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n867_), .B(new_n890_), .C1(new_n891_), .C2(new_n892_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n844_), .A2(new_n853_), .A3(new_n846_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n894_), .A2(G134gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT120), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n893_), .A2(new_n898_), .A3(new_n895_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1343gat));
  NOR4_X1   g699(.A1(new_n668_), .A2(new_n378_), .A3(new_n356_), .A4(new_n409_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n843_), .A2(new_n663_), .ZN(new_n902_));
  OAI211_X1 g701(.A(KEYINPUT121), .B(new_n901_), .C1(new_n902_), .C2(new_n806_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904_));
  INV_X1    g703(.A(new_n901_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n844_), .B2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n497_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n735_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G148gat), .ZN(G1345gat));
  AND2_X1   g710(.A1(new_n903_), .A2(new_n906_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT122), .B1(new_n912_), .B2(new_n663_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n907_), .A2(new_n914_), .A3(new_n617_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT61), .B(G155gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n913_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n916_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n914_), .B1(new_n907_), .B2(new_n617_), .ZN(new_n919_));
  AOI211_X1 g718(.A(KEYINPUT122), .B(new_n663_), .C1(new_n903_), .C2(new_n906_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n921_), .ZN(G1346gat));
  OR3_X1    g721(.A1(new_n912_), .A2(G162gat), .A3(new_n853_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G162gat), .B1(new_n912_), .B2(new_n653_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1347gat));
  NAND3_X1  g724(.A1(new_n668_), .A2(new_n409_), .A3(new_n378_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n758_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n860_), .A2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n497_), .A2(new_n265_), .ZN(new_n931_));
  XOR2_X1   g730(.A(new_n931_), .B(KEYINPUT125), .Z(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(G169gat), .B1(new_n928_), .B2(new_n498_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT62), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n935_), .A2(KEYINPUT62), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n934_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n933_), .B(new_n938_), .C1(new_n934_), .C2(new_n936_), .ZN(G1348gat));
  AOI21_X1  g738(.A(G176gat), .B1(new_n930_), .B2(new_n601_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n844_), .A2(new_n758_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n602_), .A2(new_n207_), .A3(new_n926_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(G1349gat));
  NOR2_X1   g742(.A1(new_n926_), .A2(new_n663_), .ZN(new_n944_));
  AOI21_X1  g743(.A(G183gat), .B1(new_n941_), .B2(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n663_), .A2(new_n219_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n930_), .B2(new_n946_), .ZN(G1350gat));
  NAND4_X1  g746(.A1(new_n930_), .A2(new_n260_), .A3(new_n261_), .A4(new_n661_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n930_), .A2(new_n696_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(new_n232_), .ZN(G1351gat));
  NAND3_X1  g749(.A1(new_n668_), .A2(new_n377_), .A3(new_n412_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n844_), .A2(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n497_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g753(.A1(new_n952_), .A2(new_n735_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g755(.A1(new_n844_), .A2(new_n663_), .A3(new_n951_), .ZN(new_n957_));
  AND2_X1   g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n957_), .B1(new_n958_), .B2(new_n959_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n960_), .B1(new_n957_), .B2(new_n959_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(KEYINPUT126), .ZN(G1354gat));
  AND3_X1   g761(.A1(new_n952_), .A2(G218gat), .A3(new_n696_), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n844_), .A2(new_n853_), .A3(new_n951_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n965_));
  OR2_X1    g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  AOI21_X1  g765(.A(G218gat), .B1(new_n964_), .B2(new_n965_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n963_), .B1(new_n966_), .B2(new_n967_), .ZN(G1355gat));
endmodule


