//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT85), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR3_X1   g006(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT84), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n212_));
  INV_X1    g011(.A(G141gat), .ZN(new_n213_));
  INV_X1    g012(.A(G148gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n215_), .B(new_n216_), .C1(new_n217_), .C2(new_n218_), .ZN(new_n219_));
  OAI221_X1 g018(.A(new_n205_), .B1(new_n207_), .B2(new_n208_), .C1(new_n211_), .C2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n213_), .A2(new_n214_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n207_), .A2(new_n208_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n205_), .B(KEYINPUT1), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n218_), .B(new_n221_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n225_), .A2(KEYINPUT29), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n226_), .A2(KEYINPUT28), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(KEYINPUT28), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n204_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n226_), .A2(KEYINPUT28), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n226_), .A2(KEYINPUT28), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n203_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT87), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT88), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT88), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n229_), .A2(new_n232_), .A3(new_n233_), .A4(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n229_), .A2(new_n232_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT87), .ZN(new_n240_));
  XOR2_X1   g039(.A(G211gat), .B(G218gat), .Z(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G197gat), .B(G204gat), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n241_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT21), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n241_), .A3(KEYINPUT21), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G228gat), .A2(G233gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(KEYINPUT86), .B2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(KEYINPUT29), .B2(new_n225_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(KEYINPUT86), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G78gat), .B(G106gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n254_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n256_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n240_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n238_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n258_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(new_n259_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n264_), .A2(new_n235_), .A3(new_n240_), .A4(new_n237_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G127gat), .B(G134gat), .Z(new_n268_));
  XOR2_X1   g067(.A(G113gat), .B(G120gat), .Z(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  NAND2_X1  g069(.A1(new_n225_), .A2(new_n270_), .ZN(new_n271_));
  OR3_X1    g070(.A1(new_n271_), .A2(KEYINPUT92), .A3(KEYINPUT4), .ZN(new_n272_));
  INV_X1    g071(.A(new_n225_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(KEYINPUT4), .A3(new_n271_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT92), .B1(new_n271_), .B2(KEYINPUT4), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n272_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G225gat), .A2(G233gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n275_), .A2(new_n271_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(new_n280_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G1gat), .B(G29gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G57gat), .B(G85gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT23), .ZN(new_n295_));
  OR2_X1    g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n295_), .A2(new_n296_), .B1(G169gat), .B2(G176gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT22), .B(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G169gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n301_), .B2(KEYINPUT22), .ZN(new_n302_));
  INV_X1    g101(.A(G176gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n297_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT24), .B1(new_n301_), .B2(new_n303_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  MUX2_X1   g106(.A(new_n306_), .B(KEYINPUT24), .S(new_n307_), .Z(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT26), .B(G190gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT80), .B1(new_n310_), .B2(G183gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT25), .B(G183gat), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n309_), .B(new_n311_), .C1(new_n312_), .C2(KEYINPUT80), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n308_), .A2(new_n295_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G227gat), .A2(G233gat), .ZN(new_n316_));
  INV_X1    g115(.A(G71gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(G99gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n315_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(new_n270_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G15gat), .B(G43gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT82), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT30), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT31), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n321_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n293_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n329_));
  INV_X1    g128(.A(new_n249_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(new_n305_), .A3(new_n314_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n298_), .B(KEYINPUT89), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n303_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n312_), .A2(new_n309_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n334_), .A2(new_n295_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n333_), .A2(new_n297_), .B1(new_n308_), .B2(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n331_), .B(KEYINPUT20), .C1(new_n330_), .C2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G226gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT19), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n329_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(new_n330_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n315_), .A2(new_n249_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(KEYINPUT20), .A3(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n340_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n337_), .A2(new_n329_), .A3(new_n339_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT18), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n344_), .A2(new_n352_), .A3(new_n345_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(KEYINPUT91), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT27), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT91), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n344_), .A2(new_n356_), .A3(new_n352_), .A4(new_n345_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n337_), .A2(new_n339_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n343_), .A2(new_n339_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n351_), .B(KEYINPUT27), .C1(new_n350_), .C2(new_n361_), .ZN(new_n362_));
  AND4_X1   g161(.A1(new_n267_), .A2(new_n328_), .A3(new_n358_), .A4(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n293_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n358_), .A2(new_n266_), .A3(new_n364_), .A4(new_n362_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n354_), .A2(new_n357_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n284_), .A2(new_n289_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT33), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n289_), .B1(new_n282_), .B2(new_n280_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n272_), .A2(new_n276_), .A3(new_n279_), .A4(new_n277_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT33), .B1(new_n292_), .B2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT94), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n350_), .A2(KEYINPUT32), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n361_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT94), .B1(new_n344_), .B2(new_n345_), .ZN(new_n380_));
  OAI22_X1  g179(.A1(new_n376_), .A2(new_n379_), .B1(new_n380_), .B2(new_n378_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n366_), .A2(new_n374_), .B1(new_n293_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n365_), .B1(new_n382_), .B2(new_n266_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n363_), .B1(new_n383_), .B2(new_n327_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT75), .B(G15gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G22gat), .ZN(new_n386_));
  INV_X1    g185(.A(G1gat), .ZN(new_n387_));
  INV_X1    g186(.A(G8gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT14), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G1gat), .B(G8gat), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n390_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G29gat), .B(G36gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G43gat), .B(G50gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT15), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n393_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n396_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G229gat), .A2(G233gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n396_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n401_), .B(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n406_), .B2(new_n403_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G113gat), .B(G141gat), .Z(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT79), .ZN(new_n409_));
  XOR2_X1   g208(.A(G169gat), .B(G197gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n407_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n384_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT70), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT66), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G99gat), .A2(G106gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT6), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(G99gat), .A3(G106gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT7), .ZN(new_n424_));
  INV_X1    g223(.A(G99gat), .ZN(new_n425_));
  INV_X1    g224(.A(G106gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n422_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(G85gat), .B(G92gat), .Z(new_n429_));
  AOI21_X1  g228(.A(new_n417_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT8), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n419_), .A2(new_n421_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(KEYINPUT9), .B2(new_n429_), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT10), .B(G99gat), .Z(new_n434_));
  XOR2_X1   g233(.A(KEYINPUT64), .B(G106gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT65), .B(G92gat), .ZN(new_n436_));
  INV_X1    g235(.A(G85gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n437_), .A2(KEYINPUT9), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n434_), .A2(new_n435_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n430_), .A2(new_n431_), .B1(new_n433_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n427_), .A2(new_n423_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n429_), .B1(new_n432_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT66), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n428_), .A2(new_n417_), .A3(new_n429_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(KEYINPUT8), .A3(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G57gat), .B(G64gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT11), .ZN(new_n447_));
  XOR2_X1   g246(.A(G71gat), .B(G78gat), .Z(new_n448_));
  OR2_X1    g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n446_), .A2(KEYINPUT11), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n448_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n440_), .A2(new_n445_), .A3(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n453_), .A2(KEYINPUT67), .ZN(new_n454_));
  INV_X1    g253(.A(new_n452_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n443_), .A2(KEYINPUT8), .A3(new_n444_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n433_), .A2(new_n439_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n443_), .B2(KEYINPUT8), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n455_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT68), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n452_), .B1(new_n440_), .B2(new_n445_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT68), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n453_), .A2(KEYINPUT67), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n454_), .A2(new_n460_), .A3(new_n463_), .A4(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G230gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT12), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n459_), .A2(KEYINPUT69), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT69), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT12), .B1(new_n461_), .B2(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n470_), .A2(new_n472_), .A3(new_n466_), .A4(new_n453_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G120gat), .B(G148gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT5), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G176gat), .B(G204gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  OAI21_X1  g277(.A(new_n416_), .B1(new_n474_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n468_), .A2(KEYINPUT70), .A3(new_n473_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n474_), .A2(new_n478_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(KEYINPUT71), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT71), .B1(new_n482_), .B2(new_n483_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT72), .ZN(new_n487_));
  OAI22_X1  g286(.A1(new_n485_), .A2(new_n486_), .B1(new_n487_), .B2(KEYINPUT13), .ZN(new_n488_));
  INV_X1    g287(.A(new_n486_), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n484_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n440_), .A2(new_n445_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n397_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n495_));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  OAI221_X1 g296(.A(new_n494_), .B1(KEYINPUT35), .B2(new_n497_), .C1(new_n405_), .C2(new_n493_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(KEYINPUT35), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  XNOR2_X1  g299(.A(G190gat), .B(G218gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G134gat), .B(G162gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n500_), .A2(KEYINPUT36), .A3(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(KEYINPUT36), .Z(new_n505_));
  AND2_X1   g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT74), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n510_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n507_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G127gat), .B(G155gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT16), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G183gat), .B(G211gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n452_), .B(new_n520_), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT76), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(new_n401_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n519_), .B1(new_n523_), .B2(KEYINPUT77), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n523_), .B2(new_n519_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(KEYINPUT17), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n515_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n415_), .A2(new_n492_), .A3(new_n530_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n531_), .A2(G1gat), .A3(new_n364_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n532_), .A2(KEYINPUT38), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(KEYINPUT38), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n384_), .A2(new_n507_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n529_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n492_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(new_n414_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n535_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n387_), .B1(new_n539_), .B2(new_n293_), .ZN(new_n540_));
  OR3_X1    g339(.A1(new_n533_), .A2(new_n534_), .A3(new_n540_), .ZN(G1324gat));
  NAND2_X1  g340(.A1(new_n358_), .A2(new_n362_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n388_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT39), .Z(new_n544_));
  INV_X1    g343(.A(new_n531_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n388_), .A3(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g347(.A(G15gat), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n539_), .B2(new_n326_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT41), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n545_), .A2(new_n549_), .A3(new_n326_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(G1326gat));
  INV_X1    g352(.A(G22gat), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n539_), .B2(new_n266_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT42), .Z(new_n556_));
  NAND2_X1  g355(.A1(new_n266_), .A2(new_n554_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT95), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n556_), .B1(new_n531_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT96), .ZN(G1327gat));
  INV_X1    g359(.A(KEYINPUT44), .ZN(new_n561_));
  INV_X1    g360(.A(new_n515_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n384_), .A2(KEYINPUT43), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT97), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n515_), .B1(new_n384_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n369_), .A2(new_n373_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n357_), .B2(new_n354_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n293_), .A2(new_n381_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n267_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n326_), .B1(new_n569_), .B2(new_n365_), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n570_), .A2(KEYINPUT97), .A3(new_n363_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT43), .B1(new_n565_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT98), .B(KEYINPUT43), .C1(new_n565_), .C2(new_n571_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n563_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n537_), .A2(new_n414_), .A3(new_n536_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n561_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n563_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n575_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT97), .B1(new_n570_), .B2(new_n363_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n383_), .A2(new_n327_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n363_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n564_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n582_), .A2(new_n585_), .A3(new_n515_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT98), .B1(new_n586_), .B2(KEYINPUT43), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n580_), .B1(new_n581_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(KEYINPUT44), .A3(new_n577_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n579_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G29gat), .B1(new_n590_), .B2(new_n364_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n536_), .A2(new_n508_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n415_), .A2(new_n492_), .A3(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT99), .Z(new_n594_));
  NOR2_X1   g393(.A1(new_n364_), .A2(G29gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT100), .Z(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n591_), .A2(new_n597_), .ZN(G1328gat));
  NAND3_X1  g397(.A1(new_n579_), .A2(new_n542_), .A3(new_n589_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(G36gat), .ZN(new_n600_));
  INV_X1    g399(.A(G36gat), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n594_), .A2(new_n601_), .A3(new_n542_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT45), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT45), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n594_), .A2(new_n604_), .A3(new_n601_), .A4(new_n542_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n600_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT46), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(KEYINPUT46), .A3(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1329gat));
  NAND2_X1  g410(.A1(new_n326_), .A2(G43gat), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n594_), .A2(new_n326_), .ZN(new_n613_));
  OAI22_X1  g412(.A1(new_n590_), .A2(new_n612_), .B1(G43gat), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g414(.A(G50gat), .B1(new_n594_), .B2(new_n266_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n590_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n266_), .A2(G50gat), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n616_), .B1(new_n617_), .B2(new_n618_), .ZN(G1331gat));
  NOR2_X1   g418(.A1(new_n492_), .A2(new_n413_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n535_), .A2(new_n536_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(G57gat), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n621_), .A2(new_n622_), .A3(new_n364_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n384_), .A2(new_n413_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT101), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n625_), .A2(new_n537_), .A3(new_n530_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n626_), .A2(KEYINPUT102), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(KEYINPUT102), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n293_), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n623_), .B1(new_n629_), .B2(new_n622_), .ZN(G1332gat));
  INV_X1    g429(.A(G64gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n626_), .A2(new_n631_), .A3(new_n542_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n542_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G64gat), .B1(new_n621_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT48), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(G1333gat));
  NAND3_X1  g435(.A1(new_n626_), .A2(new_n317_), .A3(new_n326_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G71gat), .B1(new_n621_), .B2(new_n327_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT49), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1334gat));
  INV_X1    g439(.A(G78gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n626_), .A2(new_n641_), .A3(new_n266_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G78gat), .B1(new_n621_), .B2(new_n267_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT50), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1335gat));
  NAND2_X1  g444(.A1(new_n592_), .A2(new_n537_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n625_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(G85gat), .B1(new_n648_), .B2(new_n293_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n620_), .A2(new_n529_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n576_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n293_), .A2(G85gat), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT103), .Z(new_n653_));
  AOI21_X1  g452(.A(new_n649_), .B1(new_n651_), .B2(new_n653_), .ZN(G1336gat));
  NAND2_X1  g453(.A1(new_n542_), .A2(new_n436_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT105), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n651_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n625_), .A2(new_n542_), .A3(new_n647_), .ZN(new_n658_));
  INV_X1    g457(.A(G92gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT104), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n658_), .A2(KEYINPUT104), .A3(new_n659_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT106), .Z(G1337gat));
  NAND3_X1  g462(.A1(new_n648_), .A2(new_n326_), .A3(new_n434_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n576_), .A2(new_n327_), .A3(new_n650_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(new_n425_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g466(.A1(new_n588_), .A2(new_n266_), .A3(new_n529_), .A4(new_n620_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G106gat), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT52), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n668_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n625_), .A2(new_n266_), .A3(new_n435_), .A4(new_n647_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT107), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n672_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT53), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT53), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n671_), .A2(new_n674_), .A3(new_n677_), .A4(new_n672_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1339gat));
  NAND3_X1  g478(.A1(new_n530_), .A2(new_n414_), .A3(new_n492_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT54), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n413_), .A2(new_n482_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n470_), .A2(new_n472_), .A3(new_n453_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(new_n467_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(new_n467_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT55), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n473_), .B(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n684_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n685_), .A2(new_n467_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT108), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n685_), .A2(new_n686_), .A3(new_n467_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n473_), .B(KEYINPUT55), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(KEYINPUT109), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n692_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT56), .B1(new_n699_), .B2(new_n478_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT56), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n480_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n692_), .B2(new_n698_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n683_), .B1(new_n700_), .B2(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n407_), .A2(new_n412_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n403_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n412_), .B1(new_n406_), .B2(new_n707_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n400_), .A2(new_n402_), .A3(new_n707_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n706_), .B(new_n712_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n507_), .B1(new_n705_), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT111), .B(KEYINPUT57), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT112), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n413_), .A2(new_n482_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n696_), .A2(KEYINPUT109), .A3(new_n697_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT109), .B1(new_n696_), .B2(new_n697_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n478_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n701_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n699_), .A2(new_n702_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n717_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n706_), .A2(new_n712_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n489_), .B2(new_n484_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n508_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n727_));
  INV_X1    g526(.A(new_n715_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n726_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n716_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(KEYINPUT57), .B(new_n508_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT116), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT116), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n714_), .A2(new_n733_), .A3(KEYINPUT57), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(KEYINPUT58), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n724_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n480_), .B1(new_n692_), .B2(new_n698_), .ZN(new_n741_));
  OAI22_X1  g540(.A1(new_n740_), .A2(new_n704_), .B1(new_n741_), .B2(KEYINPUT56), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n704_), .A2(new_n740_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n738_), .B(new_n739_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n515_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n722_), .A2(KEYINPUT113), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n704_), .A2(new_n740_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n721_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n738_), .B1(new_n748_), .B2(new_n739_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT115), .B1(new_n745_), .B2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n737_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n515_), .A4(new_n744_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n730_), .A2(new_n735_), .A3(new_n750_), .A4(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n682_), .B1(new_n755_), .B2(new_n529_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NOR4_X1   g556(.A1(new_n542_), .A2(new_n364_), .A3(new_n266_), .A4(new_n327_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT59), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n745_), .A2(new_n749_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n536_), .B1(new_n762_), .B2(new_n735_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(new_n682_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n765_));
  AND2_X1   g564(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n758_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  OAI22_X1  g566(.A1(new_n759_), .A2(new_n760_), .B1(new_n764_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G113gat), .B1(new_n768_), .B2(new_n414_), .ZN(new_n769_));
  INV_X1    g568(.A(G113gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n759_), .A2(new_n770_), .A3(new_n413_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1340gat));
  OAI21_X1  g571(.A(G120gat), .B1(new_n768_), .B2(new_n492_), .ZN(new_n773_));
  INV_X1    g572(.A(G120gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n492_), .B2(KEYINPUT60), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n759_), .B(new_n775_), .C1(KEYINPUT60), .C2(new_n774_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1341gat));
  OAI21_X1  g576(.A(G127gat), .B1(new_n768_), .B2(new_n529_), .ZN(new_n778_));
  INV_X1    g577(.A(G127gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n759_), .A2(new_n779_), .A3(new_n536_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1342gat));
  OAI21_X1  g580(.A(G134gat), .B1(new_n768_), .B2(new_n562_), .ZN(new_n782_));
  INV_X1    g581(.A(G134gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n759_), .A2(new_n783_), .A3(new_n507_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1343gat));
  NAND4_X1  g584(.A1(new_n633_), .A2(new_n293_), .A3(new_n266_), .A4(new_n327_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n756_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n413_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT118), .B(G141gat), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(G1344gat));
  NAND2_X1  g589(.A1(new_n787_), .A2(new_n537_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g591(.A1(new_n787_), .A2(new_n536_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT61), .B(G155gat), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(G1346gat));
  INV_X1    g594(.A(G162gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n787_), .A2(new_n796_), .A3(new_n507_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n756_), .A2(new_n562_), .A3(new_n786_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n796_), .ZN(G1347gat));
  NAND2_X1  g598(.A1(new_n542_), .A2(new_n328_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n266_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n763_), .B2(new_n682_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n413_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(G169gat), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(KEYINPUT119), .A3(G169gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(KEYINPUT62), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT119), .B1(new_n804_), .B2(G169gat), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT62), .ZN(new_n811_));
  INV_X1    g610(.A(new_n804_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n810_), .A2(new_n811_), .B1(new_n332_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n809_), .A2(new_n813_), .ZN(G1348gat));
  NAND2_X1  g613(.A1(new_n757_), .A2(new_n267_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n815_), .A2(KEYINPUT121), .ZN(new_n816_));
  INV_X1    g615(.A(new_n800_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(KEYINPUT121), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n492_), .A2(new_n303_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n803_), .A2(new_n537_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n303_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT120), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n824_), .A3(new_n303_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n819_), .A2(new_n820_), .B1(new_n823_), .B2(new_n825_), .ZN(G1349gat));
  NOR3_X1   g625(.A1(new_n802_), .A2(new_n312_), .A3(new_n529_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n816_), .A2(new_n536_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n828_));
  INV_X1    g627(.A(G183gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(G1350gat));
  OAI21_X1  g629(.A(G190gat), .B1(new_n802_), .B2(new_n562_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n507_), .A2(new_n309_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT122), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n802_), .B2(new_n833_), .ZN(G1351gat));
  NOR4_X1   g633(.A1(new_n633_), .A2(new_n293_), .A3(new_n267_), .A4(new_n326_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n756_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n413_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n537_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g640(.A(new_n529_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n756_), .A2(new_n836_), .A3(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT123), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n750_), .A2(new_n754_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n716_), .A2(new_n729_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n536_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n835_), .B(new_n842_), .C1(new_n850_), .C2(new_n682_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT123), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n845_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n851_), .A2(new_n854_), .A3(new_n845_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n851_), .B2(new_n845_), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n847_), .A2(new_n853_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT125), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n844_), .A2(KEYINPUT123), .A3(new_n846_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n852_), .B1(new_n851_), .B2(new_n845_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT125), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n861_), .B(new_n862_), .C1(new_n856_), .C2(new_n855_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n858_), .A2(new_n863_), .ZN(G1354gat));
  AND3_X1   g663(.A1(new_n837_), .A2(G218gat), .A3(new_n515_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n837_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n866_), .A2(KEYINPUT126), .A3(new_n508_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(G218gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT126), .B1(new_n866_), .B2(new_n508_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n865_), .B1(new_n868_), .B2(new_n869_), .ZN(G1355gat));
endmodule


