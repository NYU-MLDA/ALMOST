//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G85gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT9), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G92gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  AND2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NOR3_X1   g008(.A1(new_n208_), .A2(new_n209_), .A3(new_n205_), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT66), .B1(new_n207_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n205_), .B(G92gat), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n208_), .A2(new_n209_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n211_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT10), .B(G99gat), .Z(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT64), .B(G106gat), .Z(new_n225_));
  AOI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  INV_X1    g027(.A(G106gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n216_), .B1(new_n223_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT8), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT8), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n235_), .B(new_n216_), .C1(new_n223_), .C2(new_n232_), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n220_), .A2(new_n226_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT11), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT67), .B(G71gat), .ZN(new_n240_));
  INV_X1    g039(.A(G78gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n240_), .B(G78gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n237_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n203_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n237_), .A2(new_n247_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT68), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n248_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT12), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n237_), .B2(new_n247_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n243_), .A2(new_n246_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n234_), .A2(new_n236_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n223_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n224_), .A2(new_n225_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n211_), .B2(new_n219_), .ZN(new_n261_));
  OAI211_X1 g060(.A(KEYINPUT12), .B(new_n256_), .C1(new_n257_), .C2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n255_), .A2(new_n262_), .A3(new_n203_), .A4(new_n251_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n253_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT5), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G176gat), .B(G204gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n268_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n253_), .A2(new_n263_), .A3(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(KEYINPUT13), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT13), .B1(new_n269_), .B2(new_n271_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n202_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(KEYINPUT69), .A3(new_n272_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G225gat), .A2(G233gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n283_));
  NAND3_X1  g082(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT84), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n282_), .A2(KEYINPUT84), .A3(new_n283_), .A4(new_n284_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT82), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n284_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT1), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n287_), .A2(new_n288_), .A3(new_n293_), .A4(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT85), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n300_), .B1(new_n302_), .B2(KEYINPUT3), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(KEYINPUT86), .A3(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n300_), .B1(new_n302_), .B2(KEYINPUT86), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT3), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n298_), .B(KEYINPUT2), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n291_), .A2(new_n292_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n297_), .A2(new_n301_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G134gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G127gat), .ZN(new_n313_));
  INV_X1    g112(.A(G127gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G134gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G120gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G113gat), .ZN(new_n318_));
  INV_X1    g117(.A(G113gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G120gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n313_), .A2(new_n315_), .A3(new_n318_), .A4(new_n320_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT80), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT80), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n316_), .B2(new_n321_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n311_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n279_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n297_), .A2(new_n301_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n309_), .A2(new_n310_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n327_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n313_), .A2(new_n315_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n336_));
  AND4_X1   g135(.A1(new_n313_), .A2(new_n315_), .A3(new_n318_), .A4(new_n320_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n311_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(new_n338_), .A3(KEYINPUT4), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n331_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n335_), .A2(new_n338_), .A3(new_n279_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(new_n212_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT0), .B(G57gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(new_n341_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G197gat), .ZN(new_n350_));
  INV_X1    g149(.A(G204gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(KEYINPUT21), .A3(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G211gat), .B(G218gat), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT21), .B1(new_n352_), .B2(new_n353_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT88), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n354_), .B(new_n355_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G197gat), .B(G204gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT21), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n356_), .B1(new_n359_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n311_), .B2(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G22gat), .B(G50gat), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n364_), .B(new_n369_), .C1(new_n311_), .C2(new_n365_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n332_), .A2(new_n365_), .A3(new_n333_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n311_), .B2(new_n365_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G78gat), .B(G106gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT89), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n374_), .A2(new_n376_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n380_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n372_), .A2(new_n373_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n311_), .A2(new_n365_), .A3(new_n375_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n371_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n380_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n383_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n387_), .A2(new_n370_), .A3(new_n368_), .A4(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(G15gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(G71gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT31), .B1(new_n324_), .B2(new_n326_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n325_), .B1(new_n337_), .B2(new_n336_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT31), .ZN(new_n398_));
  INV_X1    g197(.A(new_n326_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n396_), .A2(new_n400_), .A3(new_n228_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n228_), .B1(new_n396_), .B2(new_n400_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n395_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n398_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n324_), .A2(KEYINPUT31), .A3(new_n326_), .ZN(new_n405_));
  OAI21_X1  g204(.A(G99gat), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n396_), .A2(new_n400_), .A3(new_n228_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n394_), .A3(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT79), .B(G43gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n403_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(KEYINPUT76), .A2(G169gat), .A3(G176gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n419_));
  INV_X1    g218(.A(G183gat), .ZN(new_n420_));
  INV_X1    g219(.A(G190gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n418_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G169gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT78), .B1(new_n424_), .B2(KEYINPUT22), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT22), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(G169gat), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT77), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n427_), .B2(G169gat), .ZN(new_n431_));
  INV_X1    g230(.A(G176gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n424_), .A2(KEYINPUT77), .A3(KEYINPUT22), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n416_), .B(new_n423_), .C1(new_n429_), .C2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT24), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n424_), .A2(new_n432_), .A3(KEYINPUT75), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT75), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(G169gat), .B2(G176gat), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n436_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n439_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n415_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT24), .A3(new_n413_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n440_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT26), .B1(new_n421_), .B2(KEYINPUT74), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT74), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT26), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(G190gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n420_), .A2(KEYINPUT25), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT25), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G183gat), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .A4(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n419_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(new_n417_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n435_), .B1(new_n445_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT30), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n438_), .A2(G169gat), .A3(G176gat), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT75), .B1(new_n424_), .B2(new_n432_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT24), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n414_), .A2(new_n415_), .A3(new_n436_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(new_n441_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n453_), .A2(new_n455_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(KEYINPUT30), .A3(new_n435_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n459_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT81), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT81), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n459_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n411_), .A2(new_n412_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n472_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n401_), .A2(new_n402_), .A3(new_n395_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n394_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n409_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n403_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n474_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n390_), .B1(new_n473_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n472_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n386_), .A2(new_n389_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n349_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n457_), .A2(new_n364_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n360_), .A2(new_n361_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT88), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(new_n362_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n427_), .A2(G169gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n424_), .A2(KEYINPUT22), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n432_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n423_), .A2(new_n416_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n448_), .A2(G190gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n421_), .A2(KEYINPUT26), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(new_n450_), .A3(new_n452_), .A4(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n436_), .B1(G169gat), .B2(G176gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(new_n424_), .B2(new_n432_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n455_), .B(new_n496_), .C1(new_n440_), .C2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n489_), .A2(new_n356_), .A3(new_n493_), .A4(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G226gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT19), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n486_), .A2(new_n500_), .A3(KEYINPUT20), .A4(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n504_), .A2(KEYINPUT91), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(KEYINPUT91), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n499_), .A2(new_n493_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n364_), .B2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n466_), .A2(new_n489_), .A3(new_n356_), .A4(new_n435_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n507_), .B1(new_n512_), .B2(new_n502_), .ZN(new_n513_));
  AOI211_X1 g312(.A(KEYINPUT90), .B(new_n503_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n514_));
  OAI22_X1  g313(.A1(new_n505_), .A2(new_n506_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G8gat), .B(G36gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT18), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G64gat), .B(G92gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n512_), .A2(new_n502_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT90), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n512_), .A2(new_n507_), .A3(new_n502_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n519_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n364_), .A2(new_n509_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(new_n508_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(new_n503_), .A4(new_n486_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n504_), .A2(KEYINPUT91), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(new_n525_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n520_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT93), .B(KEYINPUT27), .Z(new_n534_));
  INV_X1    g333(.A(KEYINPUT27), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n522_), .A2(new_n523_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n525_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n503_), .B1(new_n527_), .B2(new_n486_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n512_), .A2(new_n502_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n519_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT92), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT92), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n542_), .B(new_n519_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n533_), .A2(new_n534_), .B1(new_n537_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n525_), .A2(KEYINPUT32), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n524_), .A2(new_n531_), .A3(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT32), .B(new_n525_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n547_), .B(new_n548_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n335_), .A2(new_n338_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n279_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n345_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n339_), .B(new_n279_), .C1(KEYINPUT4), .C2(new_n335_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n520_), .A2(new_n532_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT33), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n346_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n340_), .A2(KEYINPUT33), .A3(new_n341_), .A4(new_n345_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n549_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n473_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n485_), .A2(new_n545_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT34), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT35), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n207_), .A2(KEYINPUT66), .A3(new_n210_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n218_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n226_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n234_), .A2(new_n236_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G29gat), .B(G36gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G43gat), .B(G50gat), .Z(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G43gat), .B(G50gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n570_), .A2(new_n571_), .A3(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT71), .B1(new_n564_), .B2(KEYINPUT35), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT15), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n575_), .A2(KEYINPUT15), .A3(new_n577_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n567_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n585_), .B(new_n584_), .C1(new_n257_), .C2(new_n261_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n567_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n579_), .A4(new_n581_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G134gat), .B(G162gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT70), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n588_), .A2(new_n591_), .A3(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n594_), .B(new_n595_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n600_), .B2(KEYINPUT72), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT72), .ZN(new_n602_));
  AOI211_X1 g401(.A(new_n602_), .B(new_n599_), .C1(new_n588_), .C2(new_n591_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT37), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT73), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n588_), .A2(new_n591_), .A3(new_n597_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n600_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n605_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NOR4_X1   g408(.A1(new_n606_), .A2(new_n600_), .A3(KEYINPUT73), .A4(KEYINPUT37), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n604_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G15gat), .B(G22gat), .ZN(new_n612_));
  INV_X1    g411(.A(G1gat), .ZN(new_n613_));
  INV_X1    g412(.A(G8gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT14), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G1gat), .B(G8gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n256_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT16), .ZN(new_n623_));
  XOR2_X1   g422(.A(G183gat), .B(G211gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT17), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n621_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT17), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n621_), .B1(new_n628_), .B2(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n611_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n618_), .B(new_n578_), .Z(new_n632_));
  NAND2_X1  g431(.A1(G229gat), .A2(G233gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n584_), .A2(new_n618_), .A3(new_n585_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n618_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n634_), .B1(new_n636_), .B2(new_n578_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n632_), .A2(new_n634_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(G113gat), .B(G141gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(G169gat), .B(G197gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n638_), .A2(new_n641_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NOR4_X1   g443(.A1(new_n278_), .A2(new_n562_), .A3(new_n631_), .A4(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n347_), .A2(new_n348_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT94), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n613_), .A3(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n649_), .B(new_n650_), .Z(new_n651_));
  NOR2_X1   g450(.A1(new_n562_), .A2(new_n607_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n652_), .A2(KEYINPUT96), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(KEYINPUT96), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n630_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n276_), .A2(new_n272_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n644_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n655_), .A2(new_n656_), .A3(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(new_n349_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n651_), .B1(new_n662_), .B2(new_n613_), .ZN(G1324gat));
  INV_X1    g462(.A(new_n545_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n645_), .A2(new_n614_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n661_), .A2(new_n664_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(G8gat), .ZN(new_n668_));
  AOI211_X1 g467(.A(KEYINPUT39), .B(new_n614_), .C1(new_n661_), .C2(new_n664_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(G1325gat));
  NOR2_X1   g471(.A1(new_n473_), .A2(new_n479_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n392_), .B1(new_n661_), .B2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(KEYINPUT97), .B(KEYINPUT41), .Z(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n645_), .A2(new_n392_), .A3(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n676_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(G1326gat));
  INV_X1    g479(.A(G22gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n482_), .B(KEYINPUT98), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n645_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n661_), .B2(new_n682_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT99), .B(KEYINPUT42), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n684_), .A2(new_n685_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(G1327gat));
  NAND2_X1  g487(.A1(new_n656_), .A2(new_n607_), .ZN(new_n689_));
  NOR4_X1   g488(.A1(new_n562_), .A2(new_n657_), .A3(new_n644_), .A4(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n349_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT43), .B1(new_n562_), .B2(new_n611_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n480_), .A2(new_n484_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n545_), .A3(new_n646_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n560_), .A2(new_n561_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  INV_X1    g496(.A(new_n611_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n696_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n692_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n660_), .A2(new_n630_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n700_), .A2(KEYINPUT44), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n648_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n691_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n713_));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n690_), .A2(new_n714_), .A3(new_n664_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT100), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT45), .ZN(new_n717_));
  OAI21_X1  g516(.A(G36gat), .B1(new_n706_), .B2(new_n545_), .ZN(new_n718_));
  AOI211_X1 g517(.A(new_n712_), .B(new_n713_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n719_));
  AND4_X1   g518(.A1(new_n710_), .A2(new_n717_), .A3(new_n711_), .A4(new_n718_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n674_), .A2(G43gat), .ZN(new_n723_));
  OR3_X1    g522(.A1(new_n706_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n706_), .B2(new_n723_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n690_), .A2(new_n674_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n724_), .B(new_n725_), .C1(G43gat), .C2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n690_), .B2(new_n682_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n482_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n707_), .B2(new_n730_), .ZN(G1331gat));
  NOR4_X1   g530(.A1(new_n562_), .A2(new_n658_), .A3(new_n631_), .A4(new_n659_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n648_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n278_), .ZN(new_n734_));
  NOR4_X1   g533(.A1(new_n655_), .A2(new_n656_), .A3(new_n659_), .A4(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT103), .B(G57gat), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n646_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n733_), .B1(new_n735_), .B2(new_n737_), .ZN(G1332gat));
  INV_X1    g537(.A(G64gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n735_), .B2(new_n664_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n732_), .A2(new_n739_), .A3(new_n664_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n735_), .B2(new_n674_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NOR2_X1   g546(.A1(new_n673_), .A2(G71gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT105), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n732_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(G1334gat));
  AOI21_X1  g550(.A(new_n241_), .B1(new_n735_), .B2(new_n682_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT50), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n732_), .A2(new_n241_), .A3(new_n682_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n562_), .A2(new_n659_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n689_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n212_), .B1(new_n758_), .B2(new_n647_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT106), .Z(new_n760_));
  NAND3_X1  g559(.A1(new_n657_), .A2(new_n656_), .A3(new_n644_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n692_), .B2(new_n699_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n646_), .A2(new_n204_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n760_), .B1(new_n762_), .B2(new_n763_), .ZN(G1336gat));
  AND2_X1   g563(.A1(new_n762_), .A2(new_n664_), .ZN(new_n765_));
  INV_X1    g564(.A(G92gat), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n664_), .A2(new_n766_), .ZN(new_n767_));
  OAI22_X1  g566(.A1(new_n765_), .A2(new_n766_), .B1(new_n758_), .B2(new_n767_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT107), .Z(G1337gat));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n756_), .A2(new_n757_), .A3(new_n224_), .A4(new_n674_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT109), .ZN(new_n772_));
  INV_X1    g571(.A(new_n761_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n697_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n774_));
  AOI211_X1 g573(.A(KEYINPUT43), .B(new_n611_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n674_), .B(new_n773_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n776_), .A2(KEYINPUT108), .A3(G99gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT108), .B1(new_n776_), .B2(G99gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n772_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(KEYINPUT51), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(KEYINPUT51), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(new_n772_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n776_), .A2(G99gat), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n776_), .A2(KEYINPUT108), .A3(G99gat), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n792_), .A2(KEYINPUT111), .A3(new_n784_), .A4(new_n772_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n787_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n770_), .B1(new_n783_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n787_), .A2(new_n793_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(KEYINPUT112), .C1(new_n782_), .C2(new_n781_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1338gat));
  NAND4_X1  g597(.A1(new_n756_), .A2(new_n757_), .A3(new_n225_), .A4(new_n482_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n762_), .A2(KEYINPUT113), .A3(new_n482_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(G106gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT113), .B1(new_n762_), .B2(new_n482_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(KEYINPUT52), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(KEYINPUT52), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n799_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT53), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n808_), .B(new_n799_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(G1339gat));
  NOR4_X1   g609(.A1(new_n698_), .A2(new_n657_), .A3(new_n656_), .A4(new_n659_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT54), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n659_), .A2(new_n271_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n203_), .A2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n255_), .A2(new_n262_), .A3(new_n251_), .A4(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(KEYINPUT115), .A2(G230gat), .A3(G233gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n817_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n255_), .A2(new_n262_), .A3(new_n251_), .A4(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n263_), .A2(KEYINPUT114), .A3(new_n814_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT114), .B1(new_n263_), .B2(new_n814_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n821_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n270_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n824_), .B2(new_n268_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n813_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n269_), .A2(new_n271_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n636_), .A2(new_n578_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n635_), .A3(new_n634_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n641_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n642_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n607_), .B1(new_n830_), .B2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT57), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n824_), .A2(new_n268_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n825_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n827_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n824_), .A2(KEYINPUT116), .A3(new_n826_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n835_), .A2(new_n271_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT58), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT117), .B1(new_n847_), .B2(new_n611_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n841_), .A2(new_n827_), .B1(new_n839_), .B2(new_n825_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n845_), .B1(new_n850_), .B2(new_n843_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n849_), .B(new_n698_), .C1(new_n851_), .C2(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(KEYINPUT58), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n838_), .B1(new_n854_), .B2(KEYINPUT118), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n848_), .A2(new_n852_), .A3(new_n856_), .A4(new_n853_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n812_), .B1(new_n858_), .B2(new_n656_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n647_), .A2(new_n664_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n390_), .A3(new_n674_), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT119), .Z(new_n863_));
  NAND3_X1  g662(.A1(new_n860_), .A2(new_n659_), .A3(new_n863_), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n837_), .B(KEYINPUT57), .Z(new_n865_));
  AOI21_X1  g664(.A(new_n630_), .B1(new_n865_), .B2(new_n854_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n812_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n868_));
  NAND2_X1  g667(.A1(new_n863_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n630_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n863_), .B1(new_n871_), .B2(new_n812_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n872_), .B2(KEYINPUT59), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n319_), .B1(new_n659_), .B2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n874_), .B2(new_n319_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n864_), .A2(new_n319_), .B1(new_n873_), .B2(new_n876_), .ZN(G1340gat));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n317_), .A2(KEYINPUT60), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n658_), .A2(KEYINPUT60), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n317_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n860_), .A2(new_n878_), .A3(new_n863_), .A4(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n881_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT122), .B1(new_n872_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  AOI211_X1 g684(.A(new_n734_), .B(new_n870_), .C1(KEYINPUT59), .C2(new_n872_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n317_), .ZN(G1341gat));
  NAND3_X1  g686(.A1(new_n860_), .A2(new_n630_), .A3(new_n863_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n630_), .A2(G127gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT123), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n888_), .A2(new_n314_), .B1(new_n873_), .B2(new_n890_), .ZN(G1342gat));
  NAND4_X1  g690(.A1(new_n860_), .A2(new_n312_), .A3(new_n607_), .A4(new_n863_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n611_), .B(new_n870_), .C1(KEYINPUT59), .C2(new_n872_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n312_), .ZN(G1343gat));
  XNOR2_X1  g693(.A(KEYINPUT124), .B(G141gat), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n484_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n860_), .A2(new_n897_), .A3(new_n861_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(new_n644_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n859_), .A2(new_n484_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n900_), .A2(new_n659_), .A3(new_n861_), .A4(new_n895_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(G1344gat));
  OAI21_X1  g701(.A(G148gat), .B1(new_n898_), .B2(new_n734_), .ZN(new_n903_));
  INV_X1    g702(.A(G148gat), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n900_), .A2(new_n904_), .A3(new_n278_), .A4(new_n861_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1345gat));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n898_), .B2(new_n656_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n907_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n900_), .A2(new_n630_), .A3(new_n861_), .A4(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1346gat));
  OAI21_X1  g710(.A(G162gat), .B1(new_n898_), .B2(new_n611_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n607_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(G162gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n900_), .A2(new_n861_), .A3(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n912_), .A2(new_n915_), .ZN(G1347gat));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  INV_X1    g716(.A(new_n682_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n648_), .A2(new_n545_), .A3(new_n673_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n918_), .B(new_n919_), .C1(new_n866_), .C2(new_n812_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n644_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n917_), .B1(new_n921_), .B2(new_n424_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n921_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n923_));
  OAI211_X1 g722(.A(KEYINPUT62), .B(G169gat), .C1(new_n920_), .C2(new_n644_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(G1348gat));
  INV_X1    g724(.A(new_n920_), .ZN(new_n926_));
  AOI21_X1  g725(.A(G176gat), .B1(new_n926_), .B2(new_n657_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n859_), .A2(new_n482_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n919_), .A2(new_n278_), .A3(G176gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n919_), .A2(new_n630_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n918_), .B(new_n932_), .C1(new_n866_), .C2(new_n812_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n859_), .A2(new_n482_), .A3(new_n931_), .ZN(new_n935_));
  AOI21_X1  g734(.A(G183gat), .B1(new_n935_), .B2(KEYINPUT125), .ZN(new_n936_));
  INV_X1    g735(.A(new_n931_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n860_), .A2(new_n390_), .A3(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n934_), .B1(new_n936_), .B2(new_n940_), .ZN(G1350gat));
  NAND4_X1  g740(.A1(new_n926_), .A2(new_n607_), .A3(new_n494_), .A4(new_n495_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n926_), .A2(new_n698_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n944_), .B2(G190gat), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n943_), .B(G190gat), .C1(new_n920_), .C2(new_n611_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n942_), .B1(new_n945_), .B2(new_n947_), .ZN(G1351gat));
  NOR2_X1   g747(.A1(new_n545_), .A2(new_n349_), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n897_), .B(new_n949_), .C1(new_n871_), .C2(new_n812_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n950_), .A2(new_n644_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(new_n350_), .ZN(G1352gat));
  NOR2_X1   g751(.A1(new_n950_), .A2(new_n734_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(new_n351_), .ZN(G1353gat));
  XOR2_X1   g753(.A(KEYINPUT63), .B(G211gat), .Z(new_n955_));
  NAND4_X1  g754(.A1(new_n900_), .A2(new_n630_), .A3(new_n949_), .A4(new_n955_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n957_), .B1(new_n950_), .B2(new_n656_), .ZN(new_n958_));
  AND2_X1   g757(.A1(new_n956_), .A2(new_n958_), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n950_), .B2(new_n611_), .ZN(new_n960_));
  OR2_X1    g759(.A1(new_n913_), .A2(G218gat), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n950_), .B2(new_n961_), .ZN(G1355gat));
endmodule


