//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_;
  XOR2_X1   g000(.A(G1gat), .B(G8gat), .Z(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT73), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208_));
  OAI211_X1 g007(.A(KEYINPUT73), .B(KEYINPUT14), .C1(new_n203_), .C2(new_n204_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT74), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n207_), .A2(new_n212_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n202_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n202_), .A3(new_n213_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(G43gat), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G29gat), .ZN(new_n221_));
  INV_X1    g020(.A(G36gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G43gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n217_), .ZN(new_n225_));
  AOI21_X1  g024(.A(G50gat), .B1(new_n220_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(new_n225_), .A3(G50gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n220_), .A2(new_n225_), .A3(G50gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(new_n226_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(KEYINPUT77), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n215_), .B(new_n216_), .C1(new_n231_), .C2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n216_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(new_n214_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n227_), .A2(KEYINPUT15), .A3(new_n228_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT15), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(new_n232_), .B2(new_n226_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n235_), .B1(new_n237_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n233_), .A2(KEYINPUT77), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n229_), .A2(new_n230_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n247_), .B(new_n248_), .C1(new_n236_), .C2(new_n214_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n235_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n245_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254_));
  INV_X1    g053(.A(G169gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G197gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n259_), .A2(KEYINPUT78), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n253_), .B(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G183gat), .A2(G190gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT23), .ZN(new_n263_));
  OR3_X1    g062(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(KEYINPUT81), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT80), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n263_), .A2(KEYINPUT81), .A3(new_n264_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT79), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT26), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n273_), .B1(new_n274_), .B2(G190gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT25), .B(G183gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G190gat), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n275_), .B(new_n276_), .C1(new_n277_), .C2(new_n273_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n266_), .A2(new_n271_), .A3(new_n272_), .A4(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n262_), .A2(KEYINPUT23), .ZN(new_n280_));
  MUX2_X1   g079(.A(new_n280_), .B(new_n263_), .S(KEYINPUT82), .Z(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(G183gat), .B2(G190gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n285_), .A2(new_n268_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n279_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G211gat), .B(G218gat), .Z(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT89), .B(G197gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G204gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n257_), .B2(G204gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n290_), .B1(new_n293_), .B2(KEYINPUT90), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n294_), .B(KEYINPUT21), .C1(KEYINPUT90), .C2(new_n293_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT91), .ZN(new_n296_));
  INV_X1    g095(.A(G204gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n298_), .B(KEYINPUT21), .C1(new_n257_), .C2(new_n297_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n299_), .B(new_n290_), .C1(new_n293_), .C2(KEYINPUT21), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n295_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n296_), .B1(new_n295_), .B2(new_n300_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n288_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT93), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n277_), .A2(new_n276_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n264_), .A2(new_n269_), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n307_), .B(KEYINPUT92), .Z(new_n308_));
  INV_X1    g107(.A(new_n267_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n281_), .B(new_n306_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n263_), .B1(G183gat), .B2(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n286_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n295_), .A2(new_n300_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(KEYINPUT93), .B(new_n288_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n305_), .A2(KEYINPUT20), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT19), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(KEYINPUT91), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n279_), .A2(new_n287_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n295_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n313_), .A2(new_n314_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(KEYINPUT20), .A3(new_n325_), .ZN(new_n326_));
  OR3_X1    g125(.A1(new_n326_), .A2(KEYINPUT97), .A3(new_n319_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT97), .B1(new_n326_), .B2(new_n319_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n320_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  AND4_X1   g134(.A1(KEYINPUT20), .A2(new_n324_), .A3(new_n319_), .A4(new_n325_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n319_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n317_), .B2(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(new_n334_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n339_), .A3(KEYINPUT27), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n338_), .A2(new_n334_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n338_), .A2(new_n334_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G113gat), .B(G120gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT85), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n345_), .A2(new_n346_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n349_), .A2(KEYINPUT85), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G155gat), .ZN(new_n352_));
  INV_X1    g151(.A(G162gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n353_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT86), .ZN(new_n358_));
  INV_X1    g157(.A(new_n355_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(KEYINPUT1), .B2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n361_), .B(KEYINPUT3), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n363_), .B(KEYINPUT2), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n355_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n369_), .B(new_n354_), .C1(new_n368_), .C2(new_n367_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n351_), .B1(new_n364_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT95), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n364_), .A2(new_n347_), .A3(new_n370_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n373_), .B(KEYINPUT4), .C1(new_n374_), .C2(new_n371_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376_));
  INV_X1    g175(.A(new_n371_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n376_), .B1(new_n377_), .B2(new_n372_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  OR3_X1    g181(.A1(new_n374_), .A2(new_n371_), .A3(new_n381_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G85gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT0), .ZN(new_n387_));
  INV_X1    g186(.A(G57gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n384_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n382_), .A2(new_n389_), .A3(new_n383_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n340_), .A2(new_n344_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n364_), .A2(new_n370_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT28), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT88), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n395_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n321_), .A2(new_n323_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n314_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(G228gat), .A3(G233gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n400_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n399_), .A2(new_n408_), .A3(new_n406_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G22gat), .B(G50gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n410_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n394_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n334_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT32), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n338_), .B2(KEYINPUT96), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n425_), .B1(new_n338_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n424_), .B1(new_n427_), .B2(new_n329_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n391_), .A2(new_n392_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n374_), .A2(new_n371_), .A3(new_n380_), .ZN(new_n431_));
  AOI211_X1 g230(.A(new_n389_), .B(new_n431_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT33), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n392_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n338_), .A2(new_n334_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n382_), .A2(KEYINPUT33), .A3(new_n389_), .A4(new_n383_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n434_), .A2(new_n339_), .A3(new_n435_), .A4(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n430_), .A2(new_n419_), .A3(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT83), .B(G15gat), .Z(new_n439_));
  NAND2_X1  g238(.A1(G227gat), .A2(G233gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(G43gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n441_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n288_), .B(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n444_), .B1(new_n446_), .B2(KEYINPUT84), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n288_), .B(KEYINPUT30), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT84), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n447_), .B(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n351_), .B(KEYINPUT31), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n421_), .A2(new_n438_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n340_), .A2(new_n344_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT98), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n419_), .A2(new_n393_), .A3(new_n453_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT98), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n340_), .A2(new_n344_), .A3(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n455_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G85gat), .B(G92gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G99gat), .A3(G106gat), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT7), .ZN(new_n470_));
  INV_X1    g269(.A(G99gat), .ZN(new_n471_));
  INV_X1    g270(.A(G106gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n464_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n477_), .B1(new_n463_), .B2(KEYINPUT64), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT10), .B(G99gat), .Z(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n472_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n466_), .A2(new_n468_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n484_), .A2(KEYINPUT9), .ZN(new_n485_));
  INV_X1    g284(.A(G85gat), .ZN(new_n486_));
  INV_X1    g285(.A(G92gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(KEYINPUT9), .A3(new_n484_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n482_), .A2(new_n483_), .A3(new_n485_), .A4(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n483_), .A2(new_n474_), .A3(new_n473_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(new_n478_), .A3(new_n464_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n480_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT65), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n480_), .A2(KEYINPUT65), .A3(new_n490_), .A4(new_n492_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n229_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n491_), .A2(new_n478_), .A3(new_n464_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n478_), .B1(new_n464_), .B2(new_n491_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n500_), .A2(new_n490_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n497_), .A2(KEYINPUT70), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G232gat), .A2(G233gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n503_), .B(KEYINPUT34), .Z(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n495_), .A2(new_n496_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n501_), .B1(new_n506_), .B2(new_n233_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT35), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n505_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n504_), .A2(KEYINPUT35), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n502_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT72), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT70), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n510_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n497_), .A2(KEYINPUT35), .A3(new_n501_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n514_), .B(new_n515_), .C1(new_n516_), .C2(new_n505_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n511_), .A2(new_n512_), .A3(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G190gat), .B(G218gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT71), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G134gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G162gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(KEYINPUT36), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n518_), .A2(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n511_), .A2(new_n512_), .A3(new_n517_), .A4(new_n523_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n511_), .A2(new_n517_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(KEYINPUT36), .A3(new_n522_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n527_), .A2(KEYINPUT37), .A3(new_n529_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G183gat), .B(G211gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(G155gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT76), .B(G127gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT17), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G71gat), .B(G78gat), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n545_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(new_n237_), .Z(new_n552_));
  OR2_X1    g351(.A1(new_n542_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(KEYINPUT17), .A3(new_n541_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n535_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n493_), .A2(KEYINPUT12), .A3(new_n549_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT66), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n493_), .A2(KEYINPUT66), .A3(KEYINPUT12), .A4(new_n549_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n549_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n559_), .A2(new_n560_), .B1(new_n506_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G230gat), .A2(G233gat), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n495_), .A2(new_n496_), .A3(new_n549_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n565_));
  OR2_X1    g364(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n506_), .A2(new_n561_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n564_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n563_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n573_), .B(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(KEYINPUT13), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(KEYINPUT13), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT69), .ZN(new_n584_));
  AND4_X1   g383(.A1(new_n261_), .A2(new_n462_), .A3(new_n556_), .A4(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n203_), .A3(new_n429_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT38), .ZN(new_n587_));
  INV_X1    g386(.A(new_n530_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n261_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n555_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n592_), .A2(KEYINPUT99), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n462_), .A2(new_n588_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(KEYINPUT99), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G1gat), .B1(new_n597_), .B2(new_n393_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n587_), .A2(new_n598_), .ZN(G1324gat));
  AND3_X1   g398(.A1(new_n340_), .A2(new_n344_), .A3(new_n459_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n459_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n594_), .A2(new_n595_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT100), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n594_), .A2(new_n606_), .A3(new_n595_), .A4(new_n603_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(G8gat), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT39), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n605_), .A2(new_n610_), .A3(new_n607_), .A4(G8gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n585_), .A2(new_n204_), .A3(new_n603_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(KEYINPUT40), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1325gat));
  INV_X1    g417(.A(G15gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n585_), .A2(new_n619_), .A3(new_n453_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G15gat), .B1(new_n597_), .B2(new_n454_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT101), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT101), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(KEYINPUT41), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT41), .B1(new_n622_), .B2(new_n623_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n620_), .B1(new_n624_), .B2(new_n625_), .ZN(G1326gat));
  NOR2_X1   g425(.A1(new_n419_), .A2(G22gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT102), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n585_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G22gat), .B1(new_n597_), .B2(new_n419_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n630_), .A2(KEYINPUT42), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(KEYINPUT42), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n629_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT103), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n635_), .B(new_n629_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(G1327gat));
  NOR2_X1   g436(.A1(new_n588_), .A2(new_n591_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n462_), .A2(new_n590_), .A3(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT104), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n221_), .A3(new_n429_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n453_), .B1(new_n394_), .B2(new_n420_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n602_), .A2(new_n458_), .B1(new_n643_), .B2(new_n438_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n644_), .B2(new_n534_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n462_), .A2(KEYINPUT43), .A3(new_n535_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n647_), .A2(KEYINPUT44), .A3(new_n590_), .A4(new_n555_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n645_), .A2(new_n590_), .A3(new_n555_), .A4(new_n646_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n652_), .A2(new_n429_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n641_), .B1(new_n653_), .B2(new_n221_), .ZN(G1328gat));
  NAND3_X1  g453(.A1(new_n640_), .A2(new_n222_), .A3(new_n603_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT45), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n648_), .A2(new_n603_), .A3(new_n651_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(G36gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n656_), .A2(KEYINPUT46), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1329gat));
  NAND3_X1  g462(.A1(new_n648_), .A2(new_n453_), .A3(new_n651_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G43gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n640_), .A2(new_n224_), .A3(new_n453_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT47), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1330gat));
  NAND3_X1  g468(.A1(new_n652_), .A2(G50gat), .A3(new_n420_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n640_), .A2(new_n420_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(G50gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n670_), .A2(KEYINPUT105), .A3(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1331gat));
  OAI21_X1  g476(.A(KEYINPUT106), .B1(new_n644_), .B2(new_n261_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n462_), .A2(new_n679_), .A3(new_n589_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n583_), .A3(new_n556_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n682_), .A2(new_n393_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n584_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n555_), .A2(new_n261_), .ZN(new_n685_));
  AND4_X1   g484(.A1(new_n462_), .A2(new_n588_), .A3(new_n684_), .A4(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n393_), .A2(new_n388_), .ZN(new_n687_));
  AOI22_X1  g486(.A1(new_n683_), .A2(new_n388_), .B1(new_n686_), .B2(new_n687_), .ZN(G1332gat));
  INV_X1    g487(.A(G64gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n686_), .B2(new_n603_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT48), .Z(new_n691_));
  NAND2_X1  g490(.A1(new_n603_), .A2(new_n689_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n682_), .B2(new_n692_), .ZN(G1333gat));
  INV_X1    g492(.A(G71gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n686_), .B2(new_n453_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT49), .Z(new_n696_));
  NAND2_X1  g495(.A1(new_n453_), .A2(new_n694_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT107), .Z(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n682_), .B2(new_n698_), .ZN(G1334gat));
  INV_X1    g498(.A(G78gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n686_), .B2(new_n420_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT50), .Z(new_n702_));
  OR2_X1    g501(.A1(new_n682_), .A2(G78gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n419_), .B2(new_n703_), .ZN(G1335gat));
  INV_X1    g503(.A(new_n638_), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n584_), .B(new_n705_), .C1(new_n678_), .C2(new_n680_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G85gat), .B1(new_n706_), .B2(new_n429_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n645_), .A2(new_n589_), .A3(new_n555_), .A4(new_n646_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n583_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n393_), .A2(new_n486_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(G1336gat));
  AOI21_X1  g511(.A(G92gat), .B1(new_n706_), .B2(new_n603_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n602_), .A2(new_n487_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n710_), .B2(new_n714_), .ZN(G1337gat));
  AOI21_X1  g514(.A(new_n705_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n716_), .A2(new_n481_), .A3(new_n453_), .A4(new_n684_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n708_), .A2(new_n709_), .A3(new_n454_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(new_n471_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT108), .B(new_n717_), .C1(new_n718_), .C2(new_n471_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(KEYINPUT51), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n719_), .B2(KEYINPUT51), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n721_), .A2(new_n724_), .A3(KEYINPUT51), .A4(new_n722_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1338gat));
  NAND2_X1  g527(.A1(new_n710_), .A2(new_n420_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n716_), .A2(new_n472_), .A3(new_n420_), .A4(new_n684_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n706_), .A2(KEYINPUT110), .A3(new_n472_), .A4(new_n420_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n708_), .A2(new_n709_), .A3(new_n419_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n472_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n730_), .A2(new_n735_), .A3(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(G1339gat));
  NAND3_X1  g540(.A1(new_n534_), .A2(new_n709_), .A3(new_n685_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT54), .Z(new_n743_));
  NAND3_X1  g542(.A1(new_n568_), .A2(new_n572_), .A3(new_n579_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n563_), .B1(new_n562_), .B2(new_n567_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n568_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n562_), .A2(KEYINPUT55), .A3(new_n563_), .A4(new_n567_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT56), .B1(new_n749_), .B2(new_n578_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n751_), .B(new_n579_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n261_), .B(new_n744_), .C1(new_n750_), .C2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n250_), .A2(new_n245_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(KEYINPUT112), .A3(new_n258_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n244_), .A2(new_n251_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n251_), .B1(new_n235_), .B2(new_n249_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(new_n259_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n756_), .A3(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n246_), .A2(new_n259_), .A3(new_n252_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n580_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n530_), .B1(new_n753_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT57), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT113), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(KEYINPUT57), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n559_), .A2(new_n560_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n567_), .A2(new_n569_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n746_), .B1(new_n771_), .B2(new_n571_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n568_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n748_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n578_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n751_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n749_), .A2(KEYINPUT56), .A3(new_n578_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n760_), .A2(new_n761_), .A3(new_n744_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT114), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n760_), .A2(new_n761_), .A3(new_n744_), .A4(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT58), .B1(new_n779_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n769_), .B1(new_n534_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n779_), .A2(KEYINPUT58), .A3(new_n784_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n784_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n790_), .A2(KEYINPUT115), .A3(new_n532_), .A4(new_n533_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n786_), .A2(new_n787_), .A3(new_n791_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n792_), .A2(KEYINPUT116), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(KEYINPUT116), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n768_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n743_), .B1(new_n795_), .B2(new_n555_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n603_), .A2(new_n393_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n420_), .A2(new_n454_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT59), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n767_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n792_), .A2(KEYINPUT117), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n765_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT117), .B1(new_n792_), .B2(new_n801_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n555_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n743_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808_));
  INV_X1    g607(.A(new_n799_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(G113gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT118), .B1(new_n589_), .B2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n800_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n796_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n813_), .A2(new_n261_), .A3(new_n814_), .A4(new_n809_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n813_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n815_), .A2(new_n811_), .B1(KEYINPUT118), .B2(new_n816_), .ZN(G1340gat));
  XNOR2_X1  g616(.A(KEYINPUT119), .B(G120gat), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n709_), .B2(KEYINPUT60), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n819_), .A2(KEYINPUT60), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n814_), .A2(new_n809_), .A3(new_n820_), .A4(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n800_), .A2(new_n810_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n825_), .A2(new_n684_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n826_), .B2(new_n819_), .ZN(G1341gat));
  OAI21_X1  g626(.A(G127gat), .B1(new_n555_), .B2(KEYINPUT121), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n825_), .B(new_n828_), .C1(KEYINPUT121), .C2(G127gat), .ZN(new_n829_));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n814_), .A2(new_n809_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n555_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n829_), .A2(new_n832_), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n831_), .B2(new_n588_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n800_), .A2(new_n810_), .A3(G134gat), .A4(new_n535_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT122), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n835_), .A2(new_n836_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1343gat));
  NOR3_X1   g640(.A1(new_n796_), .A2(new_n453_), .A3(new_n419_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n261_), .A3(new_n797_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g643(.A1(new_n842_), .A2(new_n684_), .A3(new_n797_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g645(.A1(new_n842_), .A2(new_n591_), .A3(new_n797_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT61), .B(G155gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT123), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n847_), .B(new_n849_), .Z(G1346gat));
  AND2_X1   g649(.A1(new_n842_), .A2(new_n797_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n530_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n534_), .A2(new_n353_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n852_), .A2(new_n353_), .B1(new_n851_), .B2(new_n853_), .ZN(G1347gat));
  INV_X1    g653(.A(KEYINPUT125), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n792_), .A2(new_n801_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n765_), .A3(new_n802_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n743_), .B1(new_n859_), .B2(new_n555_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n603_), .A2(new_n458_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n855_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n861_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n807_), .A2(KEYINPUT125), .A3(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n261_), .A3(new_n283_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n868_));
  NOR4_X1   g667(.A1(new_n860_), .A2(new_n868_), .A3(new_n589_), .A4(new_n861_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n861_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT124), .B1(new_n870_), .B2(new_n261_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n867_), .B1(new_n872_), .B2(G169gat), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n869_), .A2(new_n871_), .A3(KEYINPUT62), .A4(new_n255_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n866_), .B1(new_n873_), .B2(new_n874_), .ZN(G1348gat));
  NAND3_X1  g674(.A1(new_n862_), .A2(new_n583_), .A3(new_n864_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n284_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n876_), .A2(KEYINPUT126), .A3(new_n284_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n796_), .A2(new_n420_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n602_), .A2(new_n429_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n454_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n885_), .A2(new_n284_), .A3(new_n584_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n879_), .A2(new_n880_), .B1(new_n881_), .B2(new_n886_), .ZN(G1349gat));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n555_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G183gat), .B1(new_n881_), .B2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n555_), .A2(new_n276_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n865_), .B2(new_n890_), .ZN(G1350gat));
  NAND2_X1  g690(.A1(new_n865_), .A2(new_n535_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G190gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n865_), .A2(new_n277_), .A3(new_n530_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1351gat));
  NOR4_X1   g694(.A1(new_n796_), .A2(new_n453_), .A3(new_n419_), .A4(new_n883_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n261_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n684_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g699(.A(KEYINPUT63), .B(G211gat), .ZN(new_n901_));
  OR2_X1    g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n896_), .A2(new_n591_), .ZN(new_n903_));
  MUX2_X1   g702(.A(new_n901_), .B(new_n902_), .S(new_n903_), .Z(G1354gat));
  INV_X1    g703(.A(KEYINPUT127), .ZN(new_n905_));
  INV_X1    g704(.A(G218gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n534_), .A2(new_n906_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n896_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G218gat), .B1(new_n896_), .B2(new_n530_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n905_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n842_), .A2(new_n530_), .A3(new_n882_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n906_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n896_), .A2(new_n907_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n912_), .A2(KEYINPUT127), .A3(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n914_), .ZN(G1355gat));
endmodule


