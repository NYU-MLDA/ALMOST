//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n826_, new_n828_,
    new_n829_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT9), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G85gat), .A3(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT6), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n203_), .A2(new_n206_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n212_), .B(new_n213_), .C1(G99gat), .C2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(G99gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n215_), .B(new_n205_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT66), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n214_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n210_), .A3(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n221_), .A2(KEYINPUT67), .A3(new_n202_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT67), .B1(new_n221_), .B2(new_n202_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n210_), .A2(new_n217_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(new_n224_), .A3(new_n202_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n211_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G57gat), .B(G64gat), .Z(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G71gat), .B(G78gat), .ZN(new_n234_));
  OR3_X1    g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n234_), .A3(KEYINPUT11), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n229_), .A2(KEYINPUT12), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT12), .ZN(new_n240_));
  INV_X1    g039(.A(new_n211_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n214_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n219_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT6), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n209_), .B(new_n245_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n243_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n202_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n242_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n221_), .A2(KEYINPUT67), .A3(new_n202_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(KEYINPUT8), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n241_), .B1(new_n251_), .B2(new_n227_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n240_), .B1(new_n252_), .B2(new_n237_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n239_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G230gat), .A2(G233gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT64), .Z(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n237_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n251_), .A2(new_n227_), .ZN(new_n260_));
  AND4_X1   g059(.A1(KEYINPUT68), .A2(new_n260_), .A3(new_n211_), .A4(new_n237_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT68), .B1(new_n252_), .B2(new_n237_), .ZN(new_n262_));
  OAI22_X1  g061(.A1(new_n261_), .A2(new_n262_), .B1(new_n252_), .B2(new_n237_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n258_), .A2(new_n259_), .B1(new_n257_), .B2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G176gat), .B(G204gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n264_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n257_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n239_), .A2(new_n253_), .A3(new_n256_), .A4(new_n259_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n270_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n264_), .A2(new_n275_), .A3(new_n270_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n279_), .A3(KEYINPUT13), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT13), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n271_), .A2(new_n276_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(new_n278_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT78), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n286_));
  XOR2_X1   g085(.A(G29gat), .B(G36gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(G43gat), .B(G50gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G43gat), .B(G50gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(G29gat), .B(G36gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT75), .ZN(new_n294_));
  INV_X1    g093(.A(G1gat), .ZN(new_n295_));
  INV_X1    g094(.A(G8gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G15gat), .B(G22gat), .ZN(new_n300_));
  OAI211_X1 g099(.A(KEYINPUT74), .B(KEYINPUT14), .C1(new_n295_), .C2(new_n296_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G1gat), .B(G8gat), .Z(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  OAI21_X1  g103(.A(new_n286_), .B1(new_n294_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n293_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n302_), .B(new_n303_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(KEYINPUT76), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n294_), .A2(new_n304_), .A3(KEYINPUT77), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n293_), .B(KEYINPUT15), .Z(new_n319_));
  AOI22_X1  g118(.A1(new_n305_), .A2(new_n309_), .B1(new_n319_), .B2(new_n304_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n316_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n285_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT78), .B1(new_n320_), .B2(new_n316_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT79), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G113gat), .B(G141gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G169gat), .B(G197gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(KEYINPUT79), .B(new_n327_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT101), .B1(new_n284_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n284_), .A2(KEYINPUT101), .A3(new_n332_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n319_), .B1(new_n260_), .B2(new_n211_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n293_), .ZN(new_n338_));
  AOI211_X1 g137(.A(new_n241_), .B(new_n338_), .C1(new_n251_), .C2(new_n227_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT71), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G232gat), .A2(G233gat), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n341_), .B(KEYINPUT34), .Z(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT71), .B(new_n342_), .C1(new_n337_), .C2(new_n339_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n260_), .A2(new_n211_), .A3(new_n293_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n252_), .B2(new_n319_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT35), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n344_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT35), .B1(new_n344_), .B2(new_n345_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT72), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G190gat), .B(G218gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G134gat), .B(G162gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT36), .ZN(new_n356_));
  INV_X1    g155(.A(new_n345_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n342_), .B1(new_n347_), .B2(KEYINPUT71), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n348_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n344_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n352_), .A2(new_n356_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n355_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n364_), .A2(KEYINPUT36), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n369_), .A2(KEYINPUT102), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(KEYINPUT102), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n237_), .B(new_n304_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G231gat), .A2(G233gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT17), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G127gat), .B(G155gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G211gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT16), .B(G183gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  NOR3_X1   g180(.A1(new_n376_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(KEYINPUT17), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n376_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n373_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT26), .B(G190gat), .ZN(new_n387_));
  INV_X1    g186(.A(G183gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT80), .B1(new_n388_), .B2(KEYINPUT25), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT25), .B(G183gat), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n387_), .B(new_n389_), .C1(new_n390_), .C2(KEYINPUT80), .ZN(new_n391_));
  INV_X1    g190(.A(G190gat), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n388_), .A2(new_n392_), .A3(KEYINPUT23), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT23), .B1(new_n388_), .B2(new_n392_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT82), .ZN(new_n395_));
  NOR2_X1   g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n396_), .B(KEYINPUT81), .Z(new_n397_));
  INV_X1    g196(.A(KEYINPUT24), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G169gat), .A2(G176gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  OAI221_X1 g200(.A(new_n391_), .B1(new_n393_), .B2(new_n395_), .C1(new_n399_), .C2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G176gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(KEYINPUT22), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G169gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT22), .B(G169gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n403_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n408_), .B2(KEYINPUT83), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n409_), .A2(KEYINPUT84), .ZN(new_n410_));
  INV_X1    g209(.A(new_n393_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n394_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(G183gat), .B2(G190gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(KEYINPUT84), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n410_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n413_), .A2(new_n414_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n402_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G211gat), .B(G218gat), .Z(new_n420_));
  XOR2_X1   g219(.A(G197gat), .B(G204gat), .Z(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(KEYINPUT21), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT91), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(KEYINPUT91), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G197gat), .B(G204gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT90), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT21), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n423_), .B(new_n424_), .C1(new_n427_), .C2(new_n420_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n419_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n395_), .A2(new_n393_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G183gat), .A2(G190gat), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n400_), .B(new_n408_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n390_), .A2(new_n387_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n396_), .A2(KEYINPUT24), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n412_), .B(new_n433_), .C1(new_n401_), .C2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n429_), .B(KEYINPUT20), .C1(new_n428_), .C2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT19), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n419_), .A2(new_n428_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n436_), .A2(new_n428_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n443_), .A2(KEYINPUT94), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(KEYINPUT94), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n442_), .B(KEYINPUT20), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n441_), .B1(new_n446_), .B2(new_n440_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT32), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G8gat), .B(G36gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G92gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT18), .B(G64gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n450_), .B(new_n451_), .Z(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n447_), .B1(new_n448_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n437_), .A2(new_n439_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n455_), .B1(new_n446_), .B2(new_n439_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(KEYINPUT32), .A3(new_n452_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G113gat), .B(G120gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(G134gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT86), .B(G127gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT4), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G155gat), .B(G162gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(G141gat), .ZN(new_n465_));
  INV_X1    g264(.A(G148gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(KEYINPUT87), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT2), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G141gat), .A2(G148gat), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n467_), .A2(KEYINPUT3), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(KEYINPUT3), .B2(new_n467_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n469_), .A2(new_n468_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n464_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n474_), .A2(KEYINPUT1), .B1(new_n465_), .B2(new_n466_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n475_), .B(new_n469_), .C1(KEYINPUT1), .C2(new_n463_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n461_), .A2(new_n462_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n461_), .B(new_n477_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n478_), .B(new_n480_), .C1(new_n481_), .C2(new_n462_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n481_), .A2(new_n480_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G1gat), .B(G29gat), .ZN(new_n485_));
  INV_X1    g284(.A(G85gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT0), .B(G57gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n482_), .A2(new_n483_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n454_), .A2(new_n457_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT33), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n492_), .A2(KEYINPUT96), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT96), .B1(new_n492_), .B2(new_n495_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n479_), .B(new_n478_), .C1(new_n481_), .C2(new_n462_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n489_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT97), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n481_), .B(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n480_), .B2(new_n501_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n496_), .A2(new_n497_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT95), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n447_), .B2(new_n452_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n444_), .A2(new_n445_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n506_), .A2(KEYINPUT20), .A3(new_n439_), .A4(new_n442_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n453_), .B1(new_n507_), .B2(new_n441_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n447_), .A2(KEYINPUT95), .A3(new_n452_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n503_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n492_), .A2(new_n495_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n494_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n477_), .A2(KEYINPUT29), .ZN(new_n514_));
  XOR2_X1   g313(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n515_));
  XNOR2_X1  g314(.A(G22gat), .B(G50gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n514_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n477_), .A2(KEYINPUT29), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n428_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G228gat), .A2(G233gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  XNOR2_X1  g321(.A(G78gat), .B(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n518_), .B1(new_n524_), .B2(KEYINPUT93), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n522_), .A2(new_n523_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n525_), .B(new_n527_), .C1(KEYINPUT93), .C2(new_n524_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n518_), .B(KEYINPUT89), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(KEYINPUT92), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n522_), .A2(new_n531_), .A3(new_n523_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n526_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n528_), .B1(new_n529_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n461_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n419_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G15gat), .B(G43gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT31), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G71gat), .B(G99gat), .Z(new_n542_));
  NAND2_X1  g341(.A1(G227gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n538_), .A2(new_n540_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n541_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n544_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n513_), .A2(new_n535_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n534_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n533_), .A2(new_n529_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n546_), .A2(new_n547_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(new_n528_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n493_), .ZN(new_n555_));
  OR3_X1    g354(.A1(new_n509_), .A2(KEYINPUT27), .A3(new_n510_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n508_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT27), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .A4(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n549_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n336_), .A2(new_n386_), .A3(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(G1gat), .B1(new_n561_), .B2(new_n555_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n284_), .A2(new_n332_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n559_), .B2(new_n549_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n363_), .A2(new_n565_), .A3(new_n368_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT73), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n359_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT37), .B1(new_n568_), .B2(new_n367_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n567_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n571_), .A2(new_n572_), .A3(new_n385_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n564_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(new_n295_), .A3(new_n493_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT98), .Z(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n578_), .A2(KEYINPUT100), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(KEYINPUT100), .ZN(new_n580_));
  OAI221_X1 g379(.A(new_n562_), .B1(new_n576_), .B2(new_n577_), .C1(new_n579_), .C2(new_n580_), .ZN(G1324gat));
  NAND2_X1  g380(.A1(new_n556_), .A2(new_n558_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n336_), .A2(new_n386_), .A3(new_n582_), .A4(new_n560_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(G8gat), .A3(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n574_), .A2(new_n296_), .A3(new_n582_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n586_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g390(.A(new_n574_), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n592_), .A2(G15gat), .A3(new_n548_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G15gat), .B1(new_n561_), .B2(new_n548_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT104), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT41), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(KEYINPUT104), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n596_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n593_), .B1(new_n598_), .B2(new_n599_), .ZN(G1326gat));
  OR3_X1    g399(.A1(new_n592_), .A2(G22gat), .A3(new_n535_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G22gat), .B1(new_n561_), .B2(new_n535_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(KEYINPUT42), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(KEYINPUT42), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n601_), .B1(new_n603_), .B2(new_n604_), .ZN(G1327gat));
  NOR2_X1   g404(.A1(new_n369_), .A2(new_n384_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT106), .Z(new_n607_));
  AND2_X1   g406(.A1(new_n564_), .A2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(G29gat), .B1(new_n608_), .B2(new_n493_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n566_), .A2(new_n569_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT73), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n570_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n560_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT43), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n560_), .A2(new_n615_), .A3(new_n612_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n335_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n385_), .B1(new_n618_), .B2(new_n333_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(KEYINPUT44), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT44), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n619_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(KEYINPUT105), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n555_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n609_), .B1(new_n627_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g427(.A(G36gat), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n623_), .A2(new_n626_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n582_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n608_), .A2(new_n629_), .A3(new_n582_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT108), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT46), .ZN(new_n636_));
  OAI22_X1  g435(.A1(new_n631_), .A2(new_n634_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n636_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(G1329gat));
  NAND3_X1  g438(.A1(new_n630_), .A2(G43gat), .A3(new_n552_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT109), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n608_), .A2(new_n552_), .B1(KEYINPUT110), .B2(G43gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(KEYINPUT110), .B2(G43gat), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT111), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n630_), .A2(KEYINPUT109), .A3(G43gat), .A4(new_n552_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n642_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT47), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT47), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n642_), .A2(new_n646_), .A3(new_n650_), .A4(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(G1330gat));
  NAND2_X1  g451(.A1(new_n630_), .A2(new_n534_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n535_), .A2(G50gat), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n653_), .A2(G50gat), .B1(new_n608_), .B2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT112), .ZN(G1331gat));
  AOI21_X1  g455(.A(new_n332_), .B1(new_n549_), .B2(new_n559_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n284_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n386_), .ZN(new_n660_));
  INV_X1    g459(.A(G57gat), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n555_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n612_), .A2(new_n385_), .A3(new_n284_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n663_), .A2(KEYINPUT113), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(KEYINPUT113), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(new_n657_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n493_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n662_), .B1(new_n667_), .B2(new_n661_), .ZN(G1332gat));
  INV_X1    g467(.A(G64gat), .ZN(new_n669_));
  INV_X1    g468(.A(new_n660_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(new_n582_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT48), .Z(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n669_), .A3(new_n582_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1333gat));
  OAI21_X1  g473(.A(G71gat), .B1(new_n660_), .B2(new_n548_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT49), .ZN(new_n676_));
  INV_X1    g475(.A(G71gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n666_), .A2(new_n677_), .A3(new_n552_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1334gat));
  NAND2_X1  g478(.A1(new_n670_), .A2(new_n534_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G78gat), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(KEYINPUT114), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(KEYINPUT114), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT50), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(G78gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n666_), .A2(new_n686_), .A3(new_n534_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n685_), .A2(new_n687_), .A3(new_n688_), .ZN(G1335gat));
  NAND2_X1  g488(.A1(new_n659_), .A2(new_n607_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G85gat), .B1(new_n691_), .B2(new_n493_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n332_), .A2(new_n384_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n617_), .A2(new_n658_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n555_), .A2(new_n486_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(G1336gat));
  AOI21_X1  g496(.A(G92gat), .B1(new_n691_), .B2(new_n582_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n582_), .A2(G92gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n695_), .B2(new_n699_), .ZN(G1337gat));
  AOI21_X1  g499(.A(new_n215_), .B1(new_n695_), .B2(new_n552_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n552_), .A2(new_n204_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n691_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT115), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT51), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n703_), .B(new_n705_), .ZN(G1338gat));
  NAND3_X1  g505(.A1(new_n691_), .A2(new_n205_), .A3(new_n534_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G106gat), .B1(new_n694_), .B2(new_n535_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT52), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(KEYINPUT52), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI22_X1  g511(.A1(new_n329_), .A2(new_n330_), .B1(new_n264_), .B2(new_n270_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT12), .B1(new_n229_), .B2(new_n238_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n252_), .A2(new_n240_), .A3(new_n237_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n716_), .A2(KEYINPUT55), .A3(new_n256_), .A4(new_n259_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n261_), .A2(new_n262_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n257_), .B1(new_n718_), .B2(new_n254_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT55), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n273_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n717_), .A2(new_n719_), .A3(new_n721_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n722_), .A2(KEYINPUT56), .A3(new_n269_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT56), .B1(new_n722_), .B2(new_n269_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n713_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT116), .ZN(new_n726_));
  OR3_X1    g525(.A1(new_n322_), .A2(new_n323_), .A3(new_n327_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n328_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT117), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n320_), .A2(new_n317_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n729_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n277_), .A2(new_n279_), .A3(new_n727_), .A4(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT116), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n713_), .B(new_n735_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n726_), .A2(new_n734_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n369_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT57), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(KEYINPUT57), .A3(new_n369_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n722_), .A2(new_n269_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT56), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT118), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n722_), .A2(KEYINPUT56), .A3(new_n269_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n744_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n727_), .A2(new_n733_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n724_), .B2(KEYINPUT118), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(new_n274_), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT58), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n747_), .A2(new_n749_), .A3(KEYINPUT58), .A4(new_n274_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n752_), .B(new_n753_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n740_), .A2(new_n741_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n385_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n573_), .A2(new_n757_), .A3(new_n331_), .A4(new_n284_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n611_), .A2(new_n570_), .A3(new_n384_), .A4(new_n331_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT54), .B1(new_n759_), .B2(new_n658_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n756_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n553_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n582_), .A2(new_n555_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT119), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n553_), .B1(new_n756_), .B2(new_n761_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT119), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n764_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G113gat), .B1(new_n770_), .B2(new_n332_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT120), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT59), .B1(new_n762_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n765_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT120), .B1(new_n756_), .B2(new_n761_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n764_), .B(new_n767_), .C1(new_n775_), .C2(KEYINPUT59), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT121), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n774_), .A2(KEYINPUT121), .A3(new_n776_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n331_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n771_), .B1(new_n780_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g580(.A(G120gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n284_), .B2(KEYINPUT60), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(KEYINPUT60), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(KEYINPUT122), .B2(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n770_), .B(new_n785_), .C1(KEYINPUT122), .C2(new_n783_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n284_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n782_), .ZN(G1341gat));
  AND3_X1   g587(.A1(new_n774_), .A2(KEYINPUT121), .A3(new_n776_), .ZN(new_n789_));
  OAI211_X1 g588(.A(G127gat), .B(new_n384_), .C1(new_n789_), .C2(new_n777_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n385_), .B1(new_n766_), .B2(new_n769_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(G127gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(KEYINPUT123), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT123), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n791_), .B2(G127gat), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n790_), .A2(new_n794_), .A3(new_n796_), .ZN(G1342gat));
  AOI21_X1  g596(.A(G134gat), .B1(new_n770_), .B2(new_n373_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n612_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n800_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g600(.A(new_n550_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n762_), .A2(new_n802_), .A3(new_n764_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n331_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(new_n465_), .ZN(G1344gat));
  NOR2_X1   g604(.A1(new_n803_), .A2(new_n284_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(new_n466_), .ZN(G1345gat));
  NOR2_X1   g606(.A1(new_n803_), .A2(new_n385_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT61), .B(G155gat), .Z(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  OAI21_X1  g609(.A(G162gat), .B1(new_n803_), .B2(new_n799_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n372_), .A2(G162gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n803_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT124), .ZN(G1347gat));
  AOI21_X1  g613(.A(new_n493_), .B1(new_n756_), .B2(new_n761_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n815_), .A2(new_n582_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n763_), .ZN(new_n817_));
  OAI21_X1  g616(.A(G169gat), .B1(new_n817_), .B2(new_n331_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n816_), .A2(new_n332_), .A3(new_n407_), .A4(new_n763_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n822_), .B2(new_n819_), .ZN(G1348gat));
  NOR2_X1   g622(.A1(new_n817_), .A2(new_n284_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(new_n403_), .ZN(G1349gat));
  NOR2_X1   g624(.A1(new_n817_), .A2(new_n385_), .ZN(new_n826_));
  MUX2_X1   g625(.A(G183gat), .B(new_n390_), .S(new_n826_), .Z(G1350gat));
  OAI21_X1  g626(.A(G190gat), .B1(new_n817_), .B2(new_n799_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n373_), .A2(new_n387_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n817_), .B2(new_n829_), .ZN(G1351gat));
  AND2_X1   g629(.A1(new_n816_), .A2(new_n802_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n332_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n658_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT125), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(G204gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT125), .B(G204gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n834_), .B2(new_n837_), .ZN(G1353gat));
  NAND4_X1  g637(.A1(new_n815_), .A2(new_n384_), .A3(new_n802_), .A4(new_n582_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n840_));
  XOR2_X1   g639(.A(KEYINPUT63), .B(G211gat), .Z(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT126), .Z(G1354gat));
  AOI21_X1  g642(.A(G218gat), .B1(new_n831_), .B2(new_n373_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n612_), .A2(G218gat), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT127), .Z(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n831_), .B2(new_n846_), .ZN(G1355gat));
endmodule


