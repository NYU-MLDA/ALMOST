//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G85gat), .B(G92gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n204_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT10), .B(G99gat), .Z(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  AOI22_X1  g012(.A1(new_n208_), .A2(new_n209_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n205_), .A2(new_n206_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n207_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT65), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n207_), .A2(new_n214_), .A3(new_n218_), .A4(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n204_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n222_), .B(new_n223_), .C1(G99gat), .C2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n225_), .B(new_n209_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n211_), .A2(new_n213_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT67), .ZN(new_n230_));
  OR2_X1    g029(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n231_));
  NAND2_X1  g030(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n232_));
  AND4_X1   g031(.A1(new_n221_), .A2(new_n230_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n227_), .B(KEYINPUT70), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n228_), .B(KEYINPUT69), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n234_), .B1(new_n237_), .B2(new_n221_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n220_), .B1(new_n233_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G57gat), .B(G64gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G78gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n241_), .A2(new_n243_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n239_), .A2(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n220_), .B(new_n248_), .C1(new_n233_), .C2(new_n238_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n203_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n239_), .A2(new_n249_), .B1(KEYINPUT71), .B2(KEYINPUT12), .ZN(new_n253_));
  INV_X1    g052(.A(new_n250_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n203_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT72), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(new_n259_), .A3(new_n203_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n252_), .B1(new_n256_), .B2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G120gat), .B(G148gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT5), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G176gat), .B(G204gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n264_), .B(new_n265_), .Z(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT73), .B1(new_n262_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT12), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n250_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n239_), .A2(new_n249_), .A3(new_n255_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n251_), .A2(new_n259_), .A3(new_n203_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n259_), .B1(new_n251_), .B2(new_n203_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n271_), .B(new_n272_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n252_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n266_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n268_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n275_), .A2(new_n276_), .A3(new_n267_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT74), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n262_), .A2(new_n283_), .A3(new_n267_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(new_n285_), .A3(KEYINPUT13), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT13), .B1(new_n280_), .B2(new_n285_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n202_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n280_), .A2(new_n285_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT13), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(KEYINPUT75), .A3(new_n286_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G141gat), .ZN(new_n295_));
  INV_X1    g094(.A(G148gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT88), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(KEYINPUT88), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT89), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT90), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(KEYINPUT90), .A2(G155gat), .A3(G162gat), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n307_), .A2(KEYINPUT1), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT1), .B1(new_n307_), .B2(new_n308_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n304_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n301_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(new_n308_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n304_), .A2(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n297_), .A2(KEYINPUT3), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n297_), .A2(KEYINPUT3), .B1(new_n317_), .B2(new_n300_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n320_), .B(KEYINPUT91), .Z(new_n321_));
  AOI21_X1  g120(.A(new_n315_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n313_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT28), .ZN(new_n326_));
  INV_X1    g125(.A(G218gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G211gat), .ZN(new_n328_));
  INV_X1    g127(.A(G211gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(G218gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G197gat), .B(G204gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT92), .ZN(new_n335_));
  INV_X1    g134(.A(G204gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(G197gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(G197gat), .ZN(new_n338_));
  INV_X1    g137(.A(G197gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G204gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(KEYINPUT21), .B(new_n337_), .C1(new_n341_), .C2(new_n335_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT21), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n332_), .A2(new_n343_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n334_), .A2(new_n342_), .B1(new_n331_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n326_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G78gat), .B(G106gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT94), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G228gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G22gat), .B(G50gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n348_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G183gat), .ZN(new_n361_));
  INV_X1    g160(.A(G190gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(G169gat), .ZN(new_n365_));
  OR3_X1    g164(.A1(new_n365_), .A2(KEYINPUT22), .A3(G176gat), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n365_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT24), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(KEYINPUT85), .A2(G169gat), .A3(G176gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n370_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n370_), .B1(G169gat), .B2(G176gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n376_));
  INV_X1    g175(.A(G176gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n365_), .A3(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(new_n378_), .A3(new_n371_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n360_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n362_), .A2(KEYINPUT26), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n361_), .A2(KEYINPUT25), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n362_), .A2(KEYINPUT26), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n361_), .B2(KEYINPUT25), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(KEYINPUT83), .A3(G183gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n362_), .A2(KEYINPUT84), .A3(KEYINPUT26), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n386_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n369_), .B1(new_n380_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT30), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT86), .B(G43gat), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n395_), .A2(new_n396_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G227gat), .A2(G233gat), .ZN(new_n400_));
  INV_X1    g199(.A(G15gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G71gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n399_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G127gat), .B(G134gat), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n406_), .A2(KEYINPUT87), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(KEYINPUT87), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G113gat), .B(G120gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n407_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT31), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G99gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n397_), .A2(new_n398_), .A3(new_n403_), .ZN(new_n418_));
  OR3_X1    g217(.A1(new_n405_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n420_), .B(KEYINPUT99), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n414_), .B1(new_n313_), .B2(new_n322_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n319_), .A2(new_n321_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n315_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n426_), .A2(new_n413_), .A3(new_n412_), .A4(new_n312_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(new_n427_), .A3(KEYINPUT4), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n414_), .B(new_n429_), .C1(new_n313_), .C2(new_n322_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n422_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n421_), .B1(new_n423_), .B2(new_n427_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G85gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT0), .B(G57gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n437_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n417_), .B1(new_n405_), .B2(new_n418_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n419_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT104), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT19), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n360_), .A2(new_n363_), .B1(new_n367_), .B2(new_n366_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n374_), .A2(new_n360_), .A3(new_n379_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n451_), .A2(new_n383_), .A3(new_n384_), .A4(new_n385_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n449_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n448_), .B1(new_n453_), .B2(new_n345_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT97), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT96), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n374_), .A2(new_n456_), .A3(new_n360_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT24), .B1(new_n378_), .B2(new_n371_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n358_), .A2(new_n359_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT96), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT25), .B(G183gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT24), .B1(new_n365_), .B2(new_n377_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT95), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(KEYINPUT95), .B(KEYINPUT24), .C1(new_n365_), .C2(new_n377_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(new_n378_), .A3(new_n371_), .A4(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n457_), .A2(new_n460_), .A3(new_n462_), .A4(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n345_), .B1(new_n468_), .B2(new_n369_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n454_), .B1(new_n455_), .B2(new_n469_), .ZN(new_n470_));
  AOI211_X1 g269(.A(KEYINPUT97), .B(new_n345_), .C1(new_n468_), .C2(new_n369_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n447_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  AOI211_X1 g271(.A(new_n448_), .B(new_n447_), .C1(new_n346_), .C2(new_n394_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n468_), .A2(new_n369_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n345_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(G8gat), .B(G36gat), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT18), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G64gat), .B(G92gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n472_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n481_), .A2(KEYINPUT27), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n483_));
  AOI21_X1  g282(.A(new_n483_), .B1(new_n346_), .B2(new_n394_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n475_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n447_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT97), .B1(new_n474_), .B2(new_n345_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n447_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n469_), .A2(new_n455_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .A4(new_n454_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n480_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT98), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n481_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n472_), .A2(KEYINPUT98), .A3(new_n476_), .A4(new_n480_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n472_), .A2(new_n476_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n492_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT27), .ZN(new_n500_));
  AOI221_X4 g299(.A(new_n445_), .B1(new_n482_), .B2(new_n493_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n500_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n482_), .A2(new_n493_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT104), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n355_), .B(new_n444_), .C1(new_n501_), .C2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT105), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n480_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n494_), .B2(new_n481_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT27), .B1(new_n509_), .B2(new_n496_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n503_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n445_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n502_), .A2(KEYINPUT104), .A3(new_n503_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n514_), .A2(KEYINPUT105), .A3(new_n355_), .A4(new_n444_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n419_), .A2(new_n443_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n355_), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT33), .B(new_n439_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n440_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT33), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n423_), .A2(new_n427_), .A3(new_n421_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n522_), .A2(new_n437_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n428_), .A2(new_n422_), .A3(new_n430_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n521_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n519_), .B1(new_n520_), .B2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(new_n499_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n491_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT102), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT102), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n491_), .A2(new_n532_), .A3(new_n529_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n472_), .A2(new_n476_), .A3(new_n528_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT100), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n537_), .A3(new_n441_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT103), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n527_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n534_), .A2(new_n537_), .A3(KEYINPUT103), .A4(new_n441_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n518_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NOR4_X1   g341(.A1(new_n355_), .A2(new_n441_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n517_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n516_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT77), .B(G15gat), .ZN(new_n546_));
  INV_X1    g345(.A(G22gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(G1gat), .ZN(new_n549_));
  INV_X1    g348(.A(G8gat), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT14), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G1gat), .B(G8gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G29gat), .B(G36gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G43gat), .B(G50gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n554_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n557_), .B(KEYINPUT15), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(KEYINPUT81), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT81), .ZN(new_n564_));
  INV_X1    g363(.A(new_n562_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n564_), .B1(new_n554_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n560_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n554_), .A2(new_n557_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n559_), .B1(new_n568_), .B2(new_n558_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G169gat), .B(G197gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  AND2_X1   g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n570_), .A2(new_n573_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT82), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n294_), .A2(new_n545_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n557_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n239_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n239_), .A2(new_n562_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(new_n582_), .A3(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(KEYINPUT35), .A3(new_n584_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n581_), .A2(new_n588_), .A3(new_n582_), .A4(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT36), .Z(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n587_), .A2(new_n596_), .A3(new_n589_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(KEYINPUT37), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n590_), .A2(KEYINPUT76), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT76), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n587_), .A2(new_n601_), .A3(new_n589_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n602_), .A3(new_n594_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n597_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n599_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n554_), .B(new_n608_), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n248_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(G127gat), .B(G155gat), .Z(new_n612_));
  XOR2_X1   g411(.A(G183gat), .B(G211gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n614_), .B(new_n615_), .Z(new_n616_));
  INV_X1    g415(.A(KEYINPUT17), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n611_), .B1(KEYINPUT78), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n616_), .B(new_n617_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT80), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n621_), .A2(new_n622_), .B1(KEYINPUT78), .B2(new_n618_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n610_), .B(new_n623_), .C1(new_n622_), .C2(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n607_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n579_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n549_), .A3(new_n441_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n294_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n632_), .A2(new_n626_), .A3(new_n576_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n604_), .B(KEYINPUT106), .Z(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n533_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n532_), .B1(new_n491_), .B2(new_n529_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n441_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n535_), .B(KEYINPUT100), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n539_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n527_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n541_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n355_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n355_), .A2(new_n441_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n646_), .A2(new_n517_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n635_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n633_), .A2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n442_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n629_), .A2(new_n630_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n631_), .A2(new_n650_), .A3(new_n651_), .ZN(G1324gat));
  INV_X1    g451(.A(new_n514_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n628_), .A2(new_n550_), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n633_), .A2(new_n653_), .A3(new_n648_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n655_), .A2(new_n656_), .A3(G8gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n655_), .B2(G8gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g459(.A(new_n649_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n517_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G15gat), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(KEYINPUT108), .A3(G15gat), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n628_), .A2(new_n401_), .A3(new_n662_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n669_), .A3(new_n667_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n671_), .A2(new_n672_), .A3(new_n673_), .ZN(G1326gat));
  NAND2_X1  g473(.A1(new_n518_), .A2(new_n547_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT109), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n628_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n661_), .A2(new_n518_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(G22gat), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT42), .B(new_n547_), .C1(new_n661_), .C2(new_n518_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(G1327gat));
  NOR2_X1   g481(.A1(new_n604_), .A2(new_n625_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n579_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G29gat), .B1(new_n685_), .B2(new_n441_), .ZN(new_n686_));
  AOI211_X1 g485(.A(new_n625_), .B(new_n576_), .C1(new_n289_), .C2(new_n293_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n545_), .B2(new_n607_), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT43), .B(new_n606_), .C1(new_n516_), .C2(new_n544_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n647_), .B2(new_n606_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n545_), .A2(new_n688_), .A3(new_n607_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(KEYINPUT44), .A3(new_n687_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n693_), .A2(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n441_), .A2(G29gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n686_), .B1(new_n698_), .B2(new_n699_), .ZN(G1328gat));
  NOR3_X1   g499(.A1(new_n684_), .A2(G36gat), .A3(new_n514_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n693_), .A2(new_n653_), .A3(new_n697_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n704_), .A2(KEYINPUT110), .A3(G36gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT110), .B1(new_n704_), .B2(G36gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n703_), .B(KEYINPUT46), .C1(new_n705_), .C2(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1329gat));
  INV_X1    g510(.A(G43gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(new_n684_), .B2(new_n517_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n517_), .A2(new_n712_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT111), .B1(new_n698_), .B2(new_n716_), .ZN(new_n717_));
  AND4_X1   g516(.A1(KEYINPUT111), .A2(new_n693_), .A3(new_n697_), .A4(new_n716_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n715_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT47), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n715_), .B(new_n721_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n685_), .B2(new_n518_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n518_), .A2(G50gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n698_), .B2(new_n725_), .ZN(G1331gat));
  NOR3_X1   g525(.A1(new_n294_), .A2(new_n626_), .A3(new_n578_), .ZN(new_n727_));
  AND4_X1   g526(.A1(G57gat), .A2(new_n648_), .A3(new_n441_), .A4(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n576_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n294_), .A2(new_n647_), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n627_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n442_), .B1(new_n731_), .B2(KEYINPUT113), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n732_), .B1(KEYINPUT113), .B2(new_n731_), .ZN(new_n733_));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n728_), .B1(new_n733_), .B2(new_n734_), .ZN(G1332gat));
  OR3_X1    g534(.A1(new_n731_), .A2(G64gat), .A3(new_n514_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n648_), .A2(new_n727_), .A3(new_n653_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G64gat), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT48), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT48), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1333gat));
  NAND3_X1  g540(.A1(new_n648_), .A2(new_n727_), .A3(new_n662_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G71gat), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT49), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT49), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n517_), .A2(G71gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT114), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n744_), .A2(new_n745_), .B1(new_n731_), .B2(new_n747_), .ZN(G1334gat));
  OR3_X1    g547(.A1(new_n731_), .A2(G78gat), .A3(new_n355_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n648_), .A2(new_n727_), .A3(new_n518_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G78gat), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(KEYINPUT50), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(KEYINPUT50), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1335gat));
  AND2_X1   g553(.A1(new_n730_), .A2(new_n683_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G85gat), .B1(new_n755_), .B2(new_n441_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n625_), .A2(new_n729_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n632_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n689_), .A2(new_n690_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n759_), .A2(KEYINPUT115), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(KEYINPUT115), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n758_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n441_), .A2(G85gat), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT116), .Z(new_n764_));
  AOI21_X1  g563(.A(new_n756_), .B1(new_n762_), .B2(new_n764_), .ZN(G1336gat));
  INV_X1    g564(.A(G92gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n755_), .A2(new_n766_), .A3(new_n653_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n762_), .A2(new_n653_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n766_), .ZN(G1337gat));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n755_), .A2(new_n208_), .A3(new_n662_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n762_), .A2(new_n662_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n770_), .B(new_n771_), .C1(new_n772_), .C2(new_n225_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n225_), .B1(new_n762_), .B2(new_n662_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n771_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT51), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1338gat));
  NAND4_X1  g576(.A1(new_n730_), .A2(new_n209_), .A3(new_n518_), .A4(new_n683_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT117), .Z(new_n779_));
  NOR2_X1   g578(.A1(new_n758_), .A2(new_n355_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n209_), .B1(new_n780_), .B2(new_n696_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n781_), .A2(KEYINPUT52), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(KEYINPUT52), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n779_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g584(.A1(new_n607_), .A2(new_n626_), .A3(new_n578_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n287_), .A2(new_n288_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n275_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n256_), .A2(new_n261_), .A3(KEYINPUT55), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n271_), .A2(new_n251_), .A3(new_n272_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n203_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n793_), .A2(new_n794_), .A3(new_n797_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(new_n266_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(new_n266_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT56), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n563_), .A2(new_n566_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n804_), .A2(G229gat), .A3(G233gat), .A4(new_n558_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n568_), .A2(new_n558_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n573_), .B1(new_n806_), .B2(new_n559_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n574_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n801_), .A2(new_n803_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n801_), .A2(KEYINPUT58), .A3(new_n803_), .A4(new_n810_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n607_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n604_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n809_), .B1(new_n280_), .B2(new_n285_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n576_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n798_), .A2(new_n819_), .A3(new_n800_), .A4(new_n266_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n818_), .B(new_n820_), .C1(new_n799_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n817_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n802_), .B1(KEYINPUT119), .B2(KEYINPUT56), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n825_), .A2(KEYINPUT120), .A3(new_n820_), .A4(new_n818_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n816_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n815_), .B1(new_n827_), .B2(KEYINPUT57), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT122), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n830_), .B(new_n816_), .C1(new_n824_), .C2(new_n826_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n815_), .B(new_n833_), .C1(new_n827_), .C2(KEYINPUT57), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n829_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n791_), .B1(new_n835_), .B2(new_n626_), .ZN(new_n836_));
  NOR4_X1   g635(.A1(new_n653_), .A2(new_n517_), .A3(new_n518_), .A4(new_n442_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT59), .B1(new_n838_), .B2(KEYINPUT121), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(KEYINPUT121), .B2(new_n838_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n626_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n789_), .A2(new_n790_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n838_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  OAI22_X1  g643(.A1(new_n836_), .A2(new_n840_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845_), .B2(new_n577_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n844_), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n576_), .A2(G113gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(G1340gat));
  OAI21_X1  g648(.A(G120gat), .B1(new_n845_), .B2(new_n294_), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n294_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(KEYINPUT60), .B2(new_n851_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n850_), .B1(new_n847_), .B2(new_n853_), .ZN(G1341gat));
  OAI21_X1  g653(.A(G127gat), .B1(new_n845_), .B2(new_n626_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n626_), .A2(G127gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n847_), .B2(new_n856_), .ZN(G1342gat));
  OAI21_X1  g656(.A(G134gat), .B1(new_n845_), .B2(new_n606_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n634_), .A2(G134gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n847_), .B2(new_n859_), .ZN(G1343gat));
  NAND2_X1  g659(.A1(new_n842_), .A2(new_n843_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n514_), .A2(new_n517_), .A3(new_n518_), .A4(new_n441_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT123), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n861_), .A2(new_n862_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n862_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n729_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(G141gat), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n295_), .B(new_n729_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1344gat));
  OAI21_X1  g669(.A(new_n632_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G148gat), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n296_), .B(new_n632_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1345gat));
  OAI21_X1  g673(.A(new_n625_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n876_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n625_), .B(new_n878_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1346gat));
  OR2_X1    g679(.A1(new_n865_), .A2(new_n866_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n607_), .A2(G162gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT125), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n635_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n884_));
  INV_X1    g683(.A(G162gat), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n881_), .A2(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1347gat));
  NAND2_X1  g685(.A1(new_n653_), .A2(new_n444_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n518_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n831_), .B1(new_n828_), .B2(KEYINPUT122), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n625_), .B1(new_n889_), .B2(new_n834_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n729_), .B(new_n888_), .C1(new_n890_), .C2(new_n791_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT62), .B1(new_n891_), .B2(KEYINPUT22), .ZN(new_n892_));
  OAI21_X1  g691(.A(G169gat), .B1(new_n891_), .B2(KEYINPUT62), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(KEYINPUT62), .B(G169gat), .C1(new_n891_), .C2(KEYINPUT22), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1348gat));
  OAI21_X1  g695(.A(new_n888_), .B1(new_n890_), .B2(new_n791_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n897_), .A2(new_n294_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n518_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n294_), .A2(new_n377_), .A3(new_n887_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n898_), .A2(new_n377_), .B1(new_n899_), .B2(new_n900_), .ZN(G1349gat));
  NOR3_X1   g700(.A1(new_n897_), .A2(new_n626_), .A3(new_n461_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n899_), .A2(new_n625_), .A3(new_n653_), .A4(new_n444_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n361_), .B2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n897_), .B2(new_n606_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n635_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n897_), .B2(new_n906_), .ZN(G1351gat));
  NAND2_X1  g706(.A1(new_n644_), .A2(new_n517_), .ZN(new_n908_));
  XOR2_X1   g707(.A(new_n908_), .B(KEYINPUT126), .Z(new_n909_));
  NAND3_X1  g708(.A1(new_n861_), .A2(new_n653_), .A3(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n576_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n339_), .ZN(G1352gat));
  NOR2_X1   g711(.A1(new_n910_), .A2(new_n294_), .ZN(new_n913_));
  AND2_X1   g712(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n913_), .B2(new_n915_), .ZN(G1353gat));
  INV_X1    g716(.A(new_n910_), .ZN(new_n918_));
  AOI211_X1 g717(.A(KEYINPUT63), .B(G211gat), .C1(new_n918_), .C2(new_n625_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT63), .B(G211gat), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n910_), .A2(new_n626_), .A3(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1354gat));
  OAI21_X1  g721(.A(G218gat), .B1(new_n910_), .B2(new_n606_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n635_), .A2(new_n327_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n910_), .B2(new_n924_), .ZN(G1355gat));
endmodule


