//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n206_));
  INV_X1    g005(.A(G113gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G120gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT31), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n208_), .B(G120gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT31), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT85), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT30), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(G183gat), .B2(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT22), .B(G169gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(new_n226_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT84), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n222_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n222_), .A2(new_n231_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n220_), .A3(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT83), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT24), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT83), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n235_), .B(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n227_), .A2(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT26), .B(G190gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT82), .B1(new_n244_), .B2(G183gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT25), .B(G183gat), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n243_), .B(new_n245_), .C1(new_n246_), .C2(KEYINPUT82), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n234_), .A2(new_n238_), .A3(new_n242_), .A4(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT30), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n215_), .A2(new_n216_), .A3(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n218_), .A2(new_n230_), .A3(new_n248_), .A4(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n230_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n249_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n253_));
  AOI211_X1 g052(.A(KEYINPUT85), .B(KEYINPUT30), .C1(new_n211_), .C2(new_n214_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G15gat), .B(G43gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT86), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n255_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n251_), .B2(new_n255_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n205_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(new_n204_), .A3(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT87), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n266_), .B(KEYINPUT87), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G141gat), .A2(G148gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT29), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n268_), .A2(KEYINPUT88), .A3(new_n273_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT88), .B1(new_n268_), .B2(new_n273_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n275_), .B(KEYINPUT2), .Z(new_n282_));
  XOR2_X1   g081(.A(new_n276_), .B(KEYINPUT3), .Z(new_n283_));
  OAI22_X1  g082(.A1(new_n280_), .A2(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n278_), .A2(new_n279_), .A3(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT28), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT28), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G106gat), .ZN(new_n289_));
  INV_X1    g088(.A(G106gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(new_n290_), .A3(new_n287_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n293_), .A2(new_n294_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT89), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(KEYINPUT89), .A3(new_n300_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n279_), .B1(new_n278_), .B2(new_n284_), .ZN(new_n306_));
  OAI211_X1 g105(.A(G228gat), .B(G233gat), .C1(new_n305_), .C2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n306_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G228gat), .A2(G233gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n301_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G22gat), .B(G50gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(G78gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n307_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n292_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n307_), .A2(new_n310_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n312_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(new_n289_), .A3(new_n291_), .A4(new_n314_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n278_), .A2(new_n284_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n212_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n210_), .A2(new_n284_), .A3(new_n278_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(KEYINPUT4), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G225gat), .A2(G233gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT94), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT4), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(new_n329_), .A3(new_n212_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT95), .Z(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT0), .B(G57gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G85gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(G1gat), .B(G29gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n323_), .A2(new_n324_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n327_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT19), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT20), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n343_), .B1(new_n252_), .B2(new_n301_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n241_), .A2(KEYINPUT90), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n241_), .A2(KEYINPUT90), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n240_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n246_), .A2(new_n243_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n235_), .A2(new_n237_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n223_), .A4(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n234_), .B1(G183gat), .B2(G190gat), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n351_), .A2(KEYINPUT91), .A3(new_n229_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT91), .B1(new_n351_), .B2(new_n229_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n350_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n342_), .B(new_n344_), .C1(new_n354_), .C2(new_n301_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT20), .B1(new_n252_), .B2(new_n301_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n356_), .B1(new_n354_), .B2(new_n301_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n355_), .B1(new_n357_), .B2(new_n342_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G8gat), .B(G36gat), .Z(new_n359_));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT93), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n355_), .B(new_n363_), .C1(new_n357_), .C2(new_n342_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n358_), .A2(KEYINPUT93), .A3(new_n364_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n325_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n323_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n336_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT33), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n339_), .A2(new_n370_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n363_), .A2(KEYINPUT32), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n355_), .B(new_n376_), .C1(new_n357_), .C2(new_n342_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n373_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n336_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n351_), .A2(new_n229_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n305_), .A2(new_n350_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n342_), .B1(new_n381_), .B2(new_n344_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n342_), .B2(new_n357_), .ZN(new_n383_));
  OAI221_X1 g182(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .C1(new_n383_), .C2(new_n376_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n321_), .B1(new_n375_), .B2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n378_), .A2(new_n379_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n368_), .A2(new_n387_), .A3(new_n369_), .ZN(new_n388_));
  OAI211_X1 g187(.A(KEYINPUT27), .B(new_n367_), .C1(new_n383_), .C2(new_n363_), .ZN(new_n389_));
  AND4_X1   g188(.A1(new_n386_), .A2(new_n321_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n265_), .B1(new_n385_), .B2(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n262_), .A2(new_n264_), .A3(new_n386_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n321_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n388_), .A2(new_n389_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT76), .B(G22gat), .ZN(new_n397_));
  INV_X1    g196(.A(G15gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G1gat), .ZN(new_n400_));
  INV_X1    g199(.A(G8gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT14), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G1gat), .B(G8gat), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(new_n404_), .A3(new_n402_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT71), .B(G43gat), .ZN(new_n409_));
  INV_X1    g208(.A(G50gat), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n409_), .A2(new_n410_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G29gat), .B(G36gat), .ZN(new_n413_));
  OR3_X1    g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT15), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT15), .B1(new_n414_), .B2(new_n415_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n408_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT80), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n415_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n408_), .B(KEYINPUT80), .C1(new_n416_), .C2(new_n417_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(G229gat), .A2(G233gat), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n408_), .A2(new_n421_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G113gat), .B(G141gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(new_n225_), .ZN(new_n433_));
  INV_X1    g232(.A(G197gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n431_), .A2(KEYINPUT81), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n431_), .B2(KEYINPUT81), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n396_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT96), .ZN(new_n440_));
  XOR2_X1   g239(.A(G120gat), .B(G148gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(G204gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT5), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(new_n226_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT12), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT10), .B(G99gat), .Z(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n290_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G85gat), .B(G92gat), .Z(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT9), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT9), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(G85gat), .A3(G92gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n447_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT64), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT6), .ZN(new_n456_));
  AND2_X1   g255(.A1(G99gat), .A2(G106gat), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n457_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n452_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT65), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT7), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n462_), .B(new_n463_), .C1(G99gat), .C2(G106gat), .ZN(new_n464_));
  INV_X1    g263(.A(G99gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n290_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n448_), .B1(new_n460_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT8), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n468_), .B(new_n467_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT8), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n448_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n461_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT66), .B(G71gat), .ZN(new_n476_));
  INV_X1    g275(.A(G78gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G57gat), .B(G64gat), .Z(new_n479_));
  INV_X1    g278(.A(KEYINPUT11), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n480_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n445_), .B1(new_n475_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n475_), .A2(new_n485_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n447_), .A2(new_n449_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n489_));
  INV_X1    g288(.A(new_n457_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n455_), .A2(KEYINPUT6), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n453_), .A2(KEYINPUT64), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n488_), .A2(new_n489_), .A3(new_n495_), .A4(new_n451_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT68), .B1(new_n452_), .B2(new_n460_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n471_), .A2(new_n474_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n448_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n464_), .A2(new_n466_), .B1(KEYINPUT65), .B2(KEYINPUT7), .ZN(new_n502_));
  AOI211_X1 g301(.A(KEYINPUT8), .B(new_n501_), .C1(new_n495_), .C2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n473_), .B1(new_n472_), .B2(new_n448_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT67), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n498_), .B1(new_n500_), .B2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n482_), .A2(KEYINPUT12), .A3(new_n484_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n486_), .B(new_n487_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(G230gat), .A2(G233gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n487_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n475_), .A2(new_n485_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n444_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n510_), .A2(new_n513_), .A3(new_n444_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT70), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(KEYINPUT69), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n516_), .B2(KEYINPUT69), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n515_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n521_), .A2(new_n523_), .A3(KEYINPUT13), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT13), .B1(new_n521_), .B2(new_n523_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n408_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n485_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(KEYINPUT78), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G127gat), .B(G155gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G183gat), .B(G211gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n531_), .B(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n530_), .A2(new_n537_), .A3(new_n536_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT79), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G134gat), .ZN(new_n547_));
  INV_X1    g346(.A(G162gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n475_), .A2(new_n422_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n416_), .A2(new_n417_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n552_), .B1(new_n506_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n552_), .B(new_n561_), .C1(new_n506_), .C2(new_n553_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(KEYINPUT72), .A3(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(KEYINPUT72), .ZN(new_n564_));
  AOI211_X1 g363(.A(KEYINPUT73), .B(new_n551_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n564_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n551_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT73), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n549_), .A2(new_n550_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n563_), .A2(new_n564_), .A3(new_n551_), .A4(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n571_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT73), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n574_), .B1(new_n577_), .B2(new_n565_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n573_), .B(KEYINPUT75), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT74), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n578_), .B(new_n579_), .C1(new_n571_), .C2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n575_), .B1(new_n581_), .B2(KEYINPUT37), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n527_), .A2(new_n545_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n440_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n386_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n400_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT38), .ZN(new_n588_));
  INV_X1    g387(.A(new_n438_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n524_), .A2(new_n525_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n571_), .A2(new_n573_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n391_), .B2(new_n395_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(new_n543_), .A3(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G1gat), .B1(new_n594_), .B2(new_n386_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n588_), .A2(new_n595_), .ZN(G1324gat));
  OAI21_X1  g395(.A(G8gat), .B1(new_n594_), .B2(new_n394_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT39), .ZN(new_n598_));
  INV_X1    g397(.A(new_n394_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n401_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n584_), .B2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g401(.A(G15gat), .B1(new_n594_), .B2(new_n265_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT41), .Z(new_n604_));
  INV_X1    g403(.A(new_n265_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n585_), .A2(new_n398_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT97), .ZN(G1326gat));
  OAI21_X1  g407(.A(G22gat), .B1(new_n594_), .B2(new_n393_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT98), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT42), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n584_), .A2(G22gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n611_), .B1(new_n393_), .B2(new_n612_), .ZN(G1327gat));
  XNOR2_X1  g412(.A(new_n543_), .B(KEYINPUT79), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(new_n591_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n440_), .A2(new_n526_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(G29gat), .B1(new_n617_), .B2(new_n586_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n582_), .A2(KEYINPUT43), .A3(new_n396_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT43), .B1(new_n582_), .B2(new_n396_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n621_), .A2(KEYINPUT99), .A3(new_n590_), .A4(new_n545_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n581_), .A2(KEYINPUT37), .ZN(new_n623_));
  INV_X1    g422(.A(new_n575_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n396_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT43), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n582_), .A2(KEYINPUT43), .A3(new_n396_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n627_), .A2(new_n590_), .A3(new_n545_), .A4(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n622_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n622_), .A2(new_n631_), .A3(KEYINPUT100), .A4(new_n632_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n386_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n629_), .A2(new_n632_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(G29gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n618_), .B1(new_n637_), .B2(new_n640_), .ZN(G1328gat));
  INV_X1    g440(.A(G36gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n599_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n616_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT45), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n639_), .A2(new_n599_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n648_), .B2(new_n642_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n649_), .A2(KEYINPUT101), .A3(KEYINPUT46), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT46), .B1(new_n649_), .B2(KEYINPUT101), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1329gat));
  AOI21_X1  g451(.A(new_n265_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(G43gat), .A3(new_n639_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n616_), .A2(new_n265_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(G43gat), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT47), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT47), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n654_), .B(new_n658_), .C1(G43gat), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(G1330gat));
  AOI211_X1 g459(.A(new_n393_), .B(new_n638_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n321_), .A2(new_n410_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT102), .Z(new_n663_));
  OAI22_X1  g462(.A1(new_n661_), .A2(new_n410_), .B1(new_n616_), .B2(new_n663_), .ZN(G1331gat));
  NOR2_X1   g463(.A1(new_n526_), .A2(new_n438_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(new_n396_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n582_), .A2(new_n545_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G57gat), .B1(new_n669_), .B2(new_n586_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(new_n593_), .A3(new_n614_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT103), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(new_n586_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(new_n673_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g473(.A(G64gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n672_), .B2(new_n599_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT48), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n669_), .A2(new_n675_), .A3(new_n599_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1333gat));
  INV_X1    g478(.A(G71gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n672_), .B2(new_n605_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT49), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n669_), .A2(new_n680_), .A3(new_n605_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1334gat));
  AOI21_X1  g483(.A(new_n477_), .B1(new_n672_), .B2(new_n321_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT50), .Z(new_n686_));
  NAND2_X1  g485(.A1(new_n321_), .A2(new_n477_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT104), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n668_), .B2(new_n688_), .ZN(G1335gat));
  AND2_X1   g488(.A1(new_n666_), .A2(new_n615_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G85gat), .B1(new_n690_), .B2(new_n586_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n627_), .A2(new_n545_), .A3(new_n628_), .A4(new_n665_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n386_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n693_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g493(.A(G92gat), .B1(new_n690_), .B2(new_n599_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n692_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n599_), .A2(G92gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n696_), .B2(new_n697_), .ZN(G1337gat));
  NAND3_X1  g497(.A1(new_n690_), .A2(new_n446_), .A3(new_n605_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT105), .Z(new_n700_));
  OAI21_X1  g499(.A(G99gat), .B1(new_n692_), .B2(new_n265_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g502(.A(G106gat), .B1(new_n692_), .B2(new_n393_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT52), .ZN(new_n705_));
  AND4_X1   g504(.A1(new_n290_), .A2(new_n666_), .A3(new_n321_), .A4(new_n615_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT106), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT106), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT108), .ZN(new_n710_));
  XOR2_X1   g509(.A(KEYINPUT107), .B(KEYINPUT53), .Z(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n705_), .B(new_n712_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n710_), .A2(new_n711_), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n711_), .B1(new_n710_), .B2(new_n713_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1339gat));
  INV_X1    g515(.A(KEYINPUT54), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n667_), .A2(new_n717_), .A3(new_n589_), .A4(new_n526_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n623_), .A2(new_n624_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n719_), .A2(new_n526_), .A3(new_n589_), .A4(new_n614_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT54), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT55), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n508_), .A2(new_n509_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT55), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n724_), .B(new_n728_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n726_), .A2(new_n727_), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT110), .ZN(new_n731_));
  INV_X1    g530(.A(new_n444_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n726_), .A2(new_n733_), .A3(new_n727_), .A4(new_n729_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT56), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n731_), .A2(KEYINPUT56), .A3(new_n732_), .A4(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n435_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n427_), .A2(new_n430_), .A3(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n429_), .A2(new_n426_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n425_), .A2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n420_), .A2(KEYINPUT112), .A3(new_n423_), .A4(new_n424_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n742_), .B1(new_n746_), .B2(new_n426_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n516_), .B(new_n741_), .C1(new_n747_), .C2(new_n740_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n739_), .A2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(KEYINPUT114), .A2(KEYINPUT58), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n751_), .B(new_n752_), .Z(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n582_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n516_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n739_), .B2(new_n757_), .ZN(new_n758_));
  AOI211_X1 g557(.A(KEYINPUT111), .B(new_n756_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n741_), .B1(new_n747_), .B2(new_n740_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n758_), .A2(new_n759_), .A3(new_n761_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n762_), .A2(KEYINPUT57), .A3(new_n592_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n739_), .A2(new_n757_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT111), .ZN(new_n766_));
  INV_X1    g565(.A(new_n761_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n739_), .A2(new_n755_), .A3(new_n757_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n764_), .B1(new_n769_), .B2(new_n591_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n754_), .B1(new_n763_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n543_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n723_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n599_), .A2(new_n321_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n586_), .A3(new_n605_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G113gat), .B1(new_n776_), .B2(new_n438_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT57), .B1(new_n762_), .B2(new_n592_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n764_), .A3(new_n591_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n778_), .A2(new_n779_), .B1(new_n582_), .B2(new_n753_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n722_), .B1(new_n780_), .B2(new_n614_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT59), .ZN(new_n782_));
  INV_X1    g581(.A(new_n775_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT115), .B1(new_n776_), .B2(new_n782_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n722_), .B1(new_n780_), .B2(new_n543_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n783_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(KEYINPUT59), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n589_), .B(new_n785_), .C1(new_n786_), .C2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n777_), .B1(new_n791_), .B2(G113gat), .ZN(G1340gat));
  XOR2_X1   g591(.A(KEYINPUT116), .B(G120gat), .Z(new_n793_));
  AOI21_X1  g592(.A(new_n789_), .B1(new_n788_), .B2(KEYINPUT59), .ZN(new_n794_));
  AOI211_X1 g593(.A(KEYINPUT115), .B(new_n782_), .C1(new_n787_), .C2(new_n783_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n784_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n793_), .B1(new_n796_), .B2(new_n526_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n793_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n526_), .B2(KEYINPUT60), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n776_), .B(new_n799_), .C1(KEYINPUT60), .C2(new_n798_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(G1341gat));
  AOI21_X1  g600(.A(G127gat), .B1(new_n776_), .B2(new_n614_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n796_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(KEYINPUT117), .B(G127gat), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n772_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n802_), .B1(new_n803_), .B2(new_n805_), .ZN(G1342gat));
  AOI21_X1  g605(.A(G134gat), .B1(new_n776_), .B2(new_n592_), .ZN(new_n807_));
  INV_X1    g606(.A(G134gat), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n808_), .B(new_n785_), .C1(new_n786_), .C2(new_n790_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n809_), .B2(new_n582_), .ZN(G1343gat));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811_));
  NOR4_X1   g610(.A1(new_n605_), .A2(new_n599_), .A3(new_n386_), .A4(new_n393_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n773_), .B2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n787_), .A2(KEYINPUT118), .A3(new_n812_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n438_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n527_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g619(.A1(new_n816_), .A2(new_n614_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT61), .B(G155gat), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1346gat));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  AOI21_X1  g623(.A(G162gat), .B1(new_n816_), .B2(new_n592_), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n548_), .B(new_n719_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n816_), .A2(G162gat), .A3(new_n582_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n591_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n828_), .B(KEYINPUT119), .C1(G162gat), .C2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(G1347gat));
  NOR3_X1   g630(.A1(new_n265_), .A2(new_n394_), .A3(new_n586_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n781_), .A2(new_n393_), .A3(new_n832_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n833_), .A2(new_n589_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n834_), .A2(new_n835_), .A3(G169gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n834_), .B2(G169gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n833_), .B(KEYINPUT120), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n438_), .A2(new_n228_), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT121), .Z(new_n840_));
  OAI22_X1  g639(.A1(new_n836_), .A2(new_n837_), .B1(new_n838_), .B2(new_n840_), .ZN(G1348gat));
  NOR2_X1   g640(.A1(new_n773_), .A2(new_n321_), .ZN(new_n842_));
  AND4_X1   g641(.A1(G176gat), .A2(new_n842_), .A3(new_n527_), .A4(new_n832_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n833_), .B(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n527_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n843_), .B1(new_n846_), .B2(new_n226_), .ZN(G1349gat));
  AND2_X1   g646(.A1(new_n614_), .A2(new_n832_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G183gat), .B1(new_n842_), .B2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n772_), .A2(new_n246_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n845_), .B2(new_n850_), .ZN(G1350gat));
  OAI21_X1  g650(.A(G190gat), .B1(new_n838_), .B2(new_n719_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n845_), .A2(new_n592_), .A3(new_n243_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1351gat));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n605_), .A2(new_n586_), .A3(new_n394_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n787_), .A2(new_n321_), .A3(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n589_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n859_), .B2(new_n434_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(KEYINPUT122), .A3(G197gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(KEYINPUT123), .A3(new_n434_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n858_), .B2(G197gat), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n860_), .A2(new_n861_), .B1(new_n862_), .B2(new_n864_), .ZN(G1352gat));
  INV_X1    g664(.A(new_n857_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n527_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n543_), .A2(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT124), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n870_), .B1(new_n857_), .B2(new_n873_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n869_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT126), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n874_), .B(new_n876_), .ZN(G1354gat));
  NAND3_X1  g676(.A1(new_n866_), .A2(KEYINPUT127), .A3(new_n592_), .ZN(new_n878_));
  INV_X1    g677(.A(G218gat), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT127), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n857_), .B2(new_n591_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n879_), .A3(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n866_), .A2(G218gat), .A3(new_n582_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1355gat));
endmodule


