//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT83), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(KEYINPUT23), .B2(new_n205_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT84), .B(G176gat), .Z(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT22), .B(G169gat), .ZN(new_n214_));
  AOI22_X1  g013(.A1(new_n213_), .A2(new_n214_), .B1(G169gat), .B2(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NOR3_X1   g015(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(G169gat), .B2(G176gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n205_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n226_), .B1(new_n207_), .B2(new_n225_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n216_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT30), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(G43gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G227gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(G15gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n233_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n230_), .B(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(KEYINPUT31), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(KEYINPUT31), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n204_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n240_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n204_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n238_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G197gat), .B(G204gat), .Z(new_n247_));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n250_), .A2(KEYINPUT88), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n247_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n251_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(KEYINPUT88), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n247_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT89), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  OR3_X1    g057(.A1(new_n255_), .A2(KEYINPUT89), .A3(new_n257_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n252_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G228gat), .A2(G233gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  INV_X1    g062(.A(G141gat), .ZN(new_n264_));
  INV_X1    g063(.A(G148gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT1), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n263_), .B(new_n266_), .C1(new_n269_), .C2(new_n271_), .ZN(new_n272_));
  OR3_X1    g071(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n263_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n273_), .A2(new_n275_), .A3(new_n276_), .A4(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n267_), .B(KEYINPUT85), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n270_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n272_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT86), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n272_), .A2(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT86), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(KEYINPUT29), .A3(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n261_), .A2(new_n262_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n281_), .A2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(G228gat), .B(G233gat), .C1(new_n260_), .C2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G78gat), .B(G106gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n287_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n292_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n294_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n287_), .A2(new_n290_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n291_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n296_), .B1(new_n300_), .B2(new_n293_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT91), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT29), .B1(new_n283_), .B2(new_n285_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G22gat), .B(G50gat), .Z(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n304_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n302_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n306_), .A2(new_n302_), .A3(new_n307_), .ZN(new_n309_));
  OAI22_X1  g108(.A1(new_n298_), .A2(new_n301_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n297_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n309_), .A2(new_n308_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n300_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n246_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n283_), .A2(new_n243_), .A3(new_n285_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n281_), .A2(new_n204_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT95), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n317_), .A2(KEYINPUT95), .A3(new_n318_), .A4(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n204_), .A2(KEYINPUT4), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n283_), .A2(new_n285_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n318_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n317_), .A2(KEYINPUT4), .A3(new_n319_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT97), .ZN(new_n332_));
  XOR2_X1   g131(.A(G1gat), .B(G29gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT0), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT93), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G57gat), .B(G85gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT94), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n335_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n331_), .A2(new_n332_), .A3(new_n339_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n322_), .A2(new_n323_), .B1(new_n329_), .B2(new_n328_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT97), .B1(new_n341_), .B2(new_n338_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n338_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT98), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT98), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n340_), .A2(new_n342_), .A3(new_n346_), .A4(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT19), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n261_), .A2(new_n229_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n227_), .A2(new_n211_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n353_), .A2(new_n215_), .B1(new_n209_), .B2(new_n224_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT20), .B1(new_n260_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n351_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n261_), .A2(new_n229_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n260_), .A2(new_n354_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n351_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT20), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT18), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT92), .ZN(new_n364_));
  XOR2_X1   g163(.A(G64gat), .B(G92gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n356_), .A2(new_n368_), .A3(new_n360_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT27), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n359_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT20), .A4(new_n351_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n366_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n369_), .A2(new_n373_), .A3(KEYINPUT27), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n316_), .A2(new_n349_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT99), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n310_), .A2(new_n314_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n361_), .A2(new_n379_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n344_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n317_), .A2(KEYINPUT96), .A3(new_n319_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT96), .B1(new_n317_), .B2(new_n319_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n327_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n329_), .A2(new_n318_), .A3(new_n326_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n339_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n367_), .A2(new_n369_), .A3(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n343_), .A2(KEYINPUT33), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n343_), .A2(KEYINPUT33), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n378_), .B1(new_n382_), .B2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n315_), .A2(new_n375_), .A3(new_n345_), .A4(new_n347_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n377_), .B1(new_n394_), .B2(new_n246_), .ZN(new_n395_));
  AOI211_X1 g194(.A(KEYINPUT99), .B(new_n245_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n376_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(G36gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G29gat), .ZN(new_n399_));
  INV_X1    g198(.A(G29gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G36gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n401_), .A3(KEYINPUT72), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT72), .B1(new_n399_), .B2(new_n401_), .ZN(new_n404_));
  INV_X1    g203(.A(G50gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G43gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n232_), .A2(G50gat), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n406_), .A2(new_n407_), .A3(KEYINPUT73), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT73), .B1(new_n406_), .B2(new_n407_), .ZN(new_n409_));
  OAI22_X1  g208(.A1(new_n403_), .A2(new_n404_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n407_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT73), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT72), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n400_), .A2(G36gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n398_), .A2(G29gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n406_), .A2(new_n407_), .A3(KEYINPUT73), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n413_), .A2(new_n417_), .A3(new_n402_), .A4(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n410_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT15), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n410_), .A2(new_n419_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT15), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G15gat), .B(G22gat), .ZN(new_n425_));
  INV_X1    g224(.A(G1gat), .ZN(new_n426_));
  INV_X1    g225(.A(G8gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT14), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G1gat), .B(G8gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n422_), .A2(new_n424_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n431_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n420_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G229gat), .A2(G233gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n435_), .B(KEYINPUT81), .Z(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n423_), .A2(new_n431_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(G229gat), .A3(G233gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G113gat), .B(G141gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G169gat), .B(G197gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n437_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT82), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n437_), .A2(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n443_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G230gat), .ZN(new_n450_));
  INV_X1    g249(.A(G233gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT7), .ZN(new_n454_));
  INV_X1    g253(.A(G99gat), .ZN(new_n455_));
  INV_X1    g254(.A(G106gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n457_), .A2(new_n460_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G85gat), .B(G92gat), .Z(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT65), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(KEYINPUT65), .A3(new_n464_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(KEYINPUT8), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT8), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT64), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT9), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n464_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n460_), .A2(new_n461_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n472_), .A2(new_n473_), .A3(G85gat), .A4(G92gat), .ZN(new_n478_));
  OR2_X1    g277(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n456_), .A3(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .A4(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n469_), .A2(new_n471_), .A3(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G71gat), .B(G78gat), .ZN(new_n484_));
  INV_X1    g283(.A(G64gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G57gat), .ZN(new_n486_));
  INV_X1    g285(.A(G57gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G64gat), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n484_), .A2(KEYINPUT11), .A3(new_n486_), .A4(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n488_), .A3(KEYINPUT11), .ZN(new_n490_));
  AND2_X1   g289(.A1(G71gat), .A2(G78gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(G71gat), .A2(G78gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT11), .B1(new_n486_), .B2(new_n488_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n489_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT66), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT66), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n489_), .B(new_n498_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n453_), .B1(new_n483_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT68), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n468_), .A2(KEYINPUT8), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT65), .B1(new_n463_), .B2(new_n464_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n482_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n471_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n500_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT12), .ZN(new_n509_));
  INV_X1    g308(.A(new_n496_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT12), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n508_), .A2(new_n509_), .B1(new_n483_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n477_), .A2(new_n478_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n474_), .A2(new_n475_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G85gat), .B(G92gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n481_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n468_), .A2(KEYINPUT8), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n467_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n499_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT11), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n487_), .A2(G64gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n485_), .A2(G57gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n498_), .B1(new_n526_), .B2(new_n489_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n521_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n520_), .A2(new_n528_), .A3(new_n471_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(KEYINPUT68), .A3(new_n453_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n503_), .A2(new_n513_), .A3(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT67), .B1(new_n483_), .B2(new_n500_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n520_), .A2(new_n528_), .A3(new_n533_), .A4(new_n471_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n534_), .A3(new_n508_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n452_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G120gat), .B(G148gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT5), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G176gat), .B(G204gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n531_), .A2(new_n536_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT70), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n531_), .A2(new_n536_), .A3(KEYINPUT70), .A4(new_n540_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n531_), .A2(new_n536_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n540_), .B(KEYINPUT69), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT13), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(KEYINPUT71), .A3(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(KEYINPUT71), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(KEYINPUT71), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n545_), .A2(new_n548_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n397_), .A2(new_n449_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT34), .Z(new_n559_));
  INV_X1    g358(.A(KEYINPUT35), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n420_), .A2(new_n469_), .A3(new_n471_), .A4(new_n482_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT74), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n560_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n483_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n563_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n561_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n561_), .B(KEYINPUT76), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n562_), .A2(new_n564_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT75), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(KEYINPUT36), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n569_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT78), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n571_), .A2(new_n572_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n568_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n584_), .B2(new_n561_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n577_), .B(KEYINPUT36), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT77), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n580_), .B(new_n581_), .C1(new_n585_), .C2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n569_), .A2(new_n573_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n593_), .A2(new_n581_), .A3(KEYINPUT37), .A4(new_n580_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(G231gat), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(new_n451_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n433_), .A2(KEYINPUT79), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT79), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n431_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n598_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n599_), .A2(new_n601_), .A3(new_n598_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n510_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n604_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n496_), .A3(new_n602_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT16), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT80), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(KEYINPUT17), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n498_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n608_), .A2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n605_), .A2(new_n607_), .A3(new_n498_), .A4(new_n616_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n614_), .A2(new_n615_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT17), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n618_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n596_), .A2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n557_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(new_n426_), .A3(new_n348_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT38), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n593_), .A2(new_n580_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n397_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n449_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n555_), .A2(new_n631_), .A3(new_n623_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n349_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n627_), .A2(new_n634_), .ZN(G1324gat));
  XNOR2_X1  g434(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n636_));
  INV_X1    g435(.A(new_n375_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n637_), .A3(new_n632_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G8gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT39), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n625_), .A2(new_n427_), .A3(new_n637_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n639_), .A2(KEYINPUT39), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n638_), .B2(G8gat), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n641_), .B(new_n636_), .C1(new_n643_), .C2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n642_), .A2(new_n647_), .ZN(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n633_), .B2(new_n246_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n649_), .A2(KEYINPUT41), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(KEYINPUT41), .ZN(new_n651_));
  INV_X1    g450(.A(G15gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n625_), .A2(new_n652_), .A3(new_n245_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n651_), .A3(new_n653_), .ZN(G1326gat));
  OAI21_X1  g453(.A(G22gat), .B1(new_n633_), .B2(new_n378_), .ZN(new_n655_));
  XOR2_X1   g454(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n656_), .ZN(new_n658_));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n625_), .A2(new_n659_), .A3(new_n315_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n658_), .A3(new_n660_), .ZN(G1327gat));
  NAND2_X1  g460(.A1(new_n628_), .A2(new_n623_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT103), .Z(new_n663_));
  NAND2_X1  g462(.A1(new_n557_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G29gat), .B1(new_n665_), .B2(new_n348_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n556_), .A2(new_n449_), .A3(new_n623_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT102), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n397_), .A2(new_n596_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT43), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n397_), .A2(new_n671_), .A3(new_n596_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n668_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n400_), .B(new_n349_), .C1(new_n673_), .C2(KEYINPUT44), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(KEYINPUT44), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n666_), .B1(new_n674_), .B2(new_n675_), .ZN(G1328gat));
  NAND2_X1  g475(.A1(new_n673_), .A2(KEYINPUT44), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n637_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n673_), .A2(KEYINPUT44), .ZN(new_n679_));
  OAI21_X1  g478(.A(G36gat), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n557_), .A2(new_n398_), .A3(new_n637_), .A4(new_n663_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n680_), .A2(KEYINPUT46), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n375_), .B1(new_n673_), .B2(KEYINPUT44), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n398_), .B1(new_n675_), .B2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n688_), .B2(new_n683_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n685_), .A2(new_n689_), .ZN(G1329gat));
  OAI21_X1  g489(.A(new_n232_), .B1(new_n664_), .B2(new_n246_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n677_), .A2(G43gat), .A3(new_n245_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(new_n679_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT47), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n695_), .B(new_n691_), .C1(new_n692_), .C2(new_n679_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1330gat));
  OAI21_X1  g496(.A(new_n405_), .B1(new_n664_), .B2(new_n378_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n677_), .A2(G50gat), .A3(new_n315_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n679_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT105), .B(new_n698_), .C1(new_n699_), .C2(new_n679_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1331gat));
  AND3_X1   g503(.A1(new_n397_), .A2(new_n631_), .A3(new_n555_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n624_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n487_), .A3(new_n348_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n623_), .A2(new_n449_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n397_), .A2(new_n629_), .A3(new_n555_), .A4(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G57gat), .B1(new_n709_), .B2(new_n349_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1332gat));
  NAND3_X1  g510(.A1(new_n706_), .A2(new_n485_), .A3(new_n637_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G64gat), .B1(new_n709_), .B2(new_n375_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(KEYINPUT48), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(KEYINPUT48), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n712_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT106), .Z(G1333gat));
  NOR2_X1   g516(.A1(new_n246_), .A2(G71gat), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT107), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n706_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G71gat), .B1(new_n709_), .B2(new_n246_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(KEYINPUT49), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(KEYINPUT49), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT108), .Z(G1334gat));
  OAI21_X1  g524(.A(G78gat), .B1(new_n709_), .B2(new_n378_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT50), .ZN(new_n727_));
  INV_X1    g526(.A(G78gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n706_), .A2(new_n728_), .A3(new_n315_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1335gat));
  AND2_X1   g529(.A1(new_n705_), .A2(new_n663_), .ZN(new_n731_));
  INV_X1    g530(.A(G85gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n348_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n556_), .A2(new_n449_), .A3(new_n622_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n397_), .A2(new_n671_), .A3(new_n596_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n671_), .B1(new_n397_), .B2(new_n596_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(KEYINPUT109), .B(new_n734_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n349_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n733_), .B1(new_n741_), .B2(new_n732_), .ZN(G1336gat));
  AOI21_X1  g541(.A(G92gat), .B1(new_n731_), .B2(new_n637_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n739_), .A2(new_n740_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n637_), .A2(G92gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n745_), .B1(new_n746_), .B2(new_n747_), .ZN(G1337gat));
  NAND4_X1  g547(.A1(new_n731_), .A2(new_n479_), .A3(new_n480_), .A4(new_n245_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n246_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(new_n455_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT51), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n753_), .B(new_n749_), .C1(new_n750_), .C2(new_n455_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1338gat));
  NAND3_X1  g554(.A1(new_n731_), .A2(new_n456_), .A3(new_n315_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n315_), .B(new_n734_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(G106gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(G106gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT53), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n756_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1339gat));
  INV_X1    g564(.A(new_n436_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n768_));
  OR3_X1    g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n444_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n432_), .A2(new_n434_), .A3(new_n766_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n768_), .B1(new_n767_), .B2(new_n444_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n769_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n446_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n531_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n503_), .A2(new_n513_), .A3(new_n530_), .A4(KEYINPUT55), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT113), .B1(new_n513_), .B2(new_n529_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n508_), .A2(new_n509_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n483_), .A2(new_n512_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n779_), .A2(new_n529_), .A3(KEYINPUT113), .A4(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n452_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n776_), .B(new_n777_), .C1(new_n778_), .C2(new_n782_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n547_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n547_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n545_), .B(new_n774_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n543_), .A2(new_n544_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n776_), .A2(new_n777_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n782_), .A2(new_n778_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n547_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n547_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n790_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n787_), .A2(new_n788_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n774_), .A3(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n789_), .A2(new_n596_), .A3(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n449_), .B(new_n545_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n549_), .A2(new_n774_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n628_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OR2_X1    g602(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n800_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n803_), .A2(new_n804_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n623_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n590_), .A2(new_n594_), .A3(new_n631_), .A4(new_n622_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n555_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n809_), .A2(new_n810_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT112), .B(new_n811_), .C1(new_n555_), .C2(new_n812_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n816_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n817_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n595_), .A2(new_n551_), .A3(new_n554_), .A4(new_n708_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT112), .B1(new_n821_), .B2(new_n811_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n819_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n808_), .A2(new_n818_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n349_), .A2(new_n637_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n316_), .A4(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n316_), .A2(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n823_), .A2(new_n818_), .ZN(new_n831_));
  AOI211_X1 g630(.A(new_n773_), .B(new_n790_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n595_), .B1(new_n832_), .B2(new_n798_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n833_), .A2(new_n789_), .B1(new_n804_), .B2(new_n803_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n807_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n622_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT117), .B1(new_n831_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n808_), .A2(new_n838_), .A3(new_n818_), .A4(new_n823_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n830_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT59), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n829_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n631_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n631_), .A2(G113gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n841_), .B2(new_n845_), .ZN(G1340gat));
  OAI21_X1  g645(.A(G120gat), .B1(new_n843_), .B2(new_n556_), .ZN(new_n847_));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n556_), .B2(KEYINPUT60), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n849_), .A2(KEYINPUT119), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(KEYINPUT119), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n850_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n848_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n847_), .B1(new_n841_), .B2(new_n852_), .ZN(G1341gat));
  OAI21_X1  g652(.A(G127gat), .B1(new_n843_), .B2(new_n623_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n623_), .A2(G127gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n841_), .B2(new_n855_), .ZN(G1342gat));
  XOR2_X1   g655(.A(KEYINPUT121), .B(G134gat), .Z(new_n857_));
  NAND4_X1  g656(.A1(new_n829_), .A2(new_n842_), .A3(new_n596_), .A4(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G134gat), .B1(new_n840_), .B2(new_n628_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT120), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n859_), .A2(KEYINPUT120), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n858_), .A2(new_n860_), .A3(new_n861_), .ZN(G1343gat));
  INV_X1    g661(.A(new_n826_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n245_), .A2(new_n378_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI211_X1 g664(.A(new_n863_), .B(new_n865_), .C1(new_n837_), .C2(new_n839_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n449_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n555_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G148gat), .ZN(G1345gat));
  XOR2_X1   g669(.A(KEYINPUT61), .B(G155gat), .Z(new_n871_));
  NAND2_X1  g670(.A1(new_n837_), .A2(new_n839_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n872_), .A2(new_n622_), .A3(new_n826_), .A4(new_n864_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n865_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n877_), .A2(KEYINPUT122), .A3(new_n622_), .A4(new_n826_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n875_), .A2(new_n876_), .A3(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n876_), .B1(new_n875_), .B2(new_n878_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n871_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT122), .B1(new_n866_), .B2(new_n622_), .ZN(new_n882_));
  AND4_X1   g681(.A1(KEYINPUT122), .A2(new_n877_), .A3(new_n622_), .A4(new_n826_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT123), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n875_), .A2(new_n876_), .A3(new_n878_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n871_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n881_), .A2(new_n887_), .ZN(G1346gat));
  NAND2_X1  g687(.A1(new_n866_), .A2(new_n628_), .ZN(new_n889_));
  INV_X1    g688(.A(G162gat), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n595_), .A2(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT124), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n889_), .A2(new_n890_), .B1(new_n866_), .B2(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT125), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n348_), .A2(new_n375_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n316_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n824_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n449_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n900_));
  INV_X1    g699(.A(new_n214_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(new_n902_));
  AOI21_X1  g701(.A(KEYINPUT62), .B1(new_n899_), .B2(G169gat), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1348gat));
  AOI21_X1  g703(.A(new_n896_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(G176gat), .A3(new_n555_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n907_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n898_), .A2(new_n555_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n908_), .A2(new_n909_), .B1(new_n213_), .B2(new_n910_), .ZN(G1349gat));
  INV_X1    g710(.A(new_n898_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n912_), .A2(new_n218_), .A3(new_n623_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G183gat), .B1(new_n905_), .B2(new_n622_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n912_), .B2(new_n595_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n898_), .A2(new_n628_), .A3(new_n219_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1351gat));
  NAND3_X1  g717(.A1(new_n877_), .A2(new_n449_), .A3(new_n895_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g719(.A1(new_n877_), .A2(new_n555_), .A3(new_n895_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g721(.A(new_n623_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n877_), .A2(new_n895_), .A3(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT127), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n924_), .B(new_n926_), .Z(G1354gat));
  NAND3_X1  g726(.A1(new_n877_), .A2(new_n596_), .A3(new_n895_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(G218gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n629_), .A2(G218gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n877_), .A2(new_n895_), .A3(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1355gat));
endmodule


