//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_;
  XNOR2_X1  g000(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(KEYINPUT24), .A3(new_n206_), .ZN(new_n207_));
  OR3_X1    g006(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT25), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G183gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G190gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT26), .B1(new_n212_), .B2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n209_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT80), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n223_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n229_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n222_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT23), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT81), .B1(new_n230_), .B2(new_n228_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n214_), .A2(new_n220_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT81), .A4(KEYINPUT23), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G169gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n232_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT90), .ZN(new_n244_));
  INV_X1    g043(.A(G197gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT89), .B1(new_n245_), .B2(G204gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT89), .ZN(new_n247_));
  INV_X1    g046(.A(G204gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(G197gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(G204gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n243_), .A2(KEYINPUT90), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n244_), .A2(KEYINPUT21), .A3(new_n251_), .A4(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT21), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n246_), .A2(new_n249_), .A3(new_n254_), .A4(new_n250_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n250_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n245_), .A2(G204gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT21), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n243_), .A2(KEYINPUT90), .ZN(new_n259_));
  INV_X1    g058(.A(G218gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(G211gat), .ZN(new_n261_));
  INV_X1    g060(.A(G211gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(G218gat), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n261_), .A2(new_n263_), .A3(KEYINPUT90), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n255_), .B(new_n258_), .C1(new_n259_), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n253_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n202_), .B1(new_n242_), .B2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n253_), .A2(new_n265_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n231_), .A2(new_n236_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n240_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n235_), .A2(new_n208_), .A3(new_n237_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT93), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT93), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n235_), .A2(new_n274_), .A3(new_n208_), .A4(new_n237_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT92), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n220_), .A2(KEYINPUT26), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n211_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n276_), .B(new_n207_), .C1(new_n218_), .C2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n207_), .B1(new_n218_), .B2(new_n278_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT92), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n275_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n268_), .B(new_n270_), .C1(new_n273_), .C2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n267_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G226gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT19), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n270_), .B1(new_n273_), .B2(new_n282_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n266_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n286_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT20), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n231_), .A2(new_n222_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(new_n268_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n289_), .A2(new_n290_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n287_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT18), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n272_), .A2(new_n275_), .A3(new_n279_), .A4(new_n281_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n268_), .B1(new_n301_), .B2(new_n270_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT20), .B1(new_n242_), .B2(new_n266_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n286_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n299_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n242_), .A2(new_n266_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n283_), .A2(KEYINPUT20), .A3(new_n290_), .A4(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n300_), .A2(KEYINPUT27), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n304_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n305_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G22gat), .B(G50gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G155gat), .B(G162gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT86), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT86), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n321_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324_));
  INV_X1    g123(.A(G141gat), .ZN(new_n325_));
  INV_X1    g124(.A(G148gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT2), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n318_), .B1(new_n323_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n325_), .A2(new_n326_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n334_), .A2(new_n328_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n335_), .B(new_n336_), .C1(KEYINPUT1), .C2(new_n317_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT28), .B1(new_n338_), .B2(KEYINPUT29), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n333_), .A2(new_n340_), .A3(new_n341_), .A4(new_n337_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n316_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n338_), .A2(KEYINPUT29), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT88), .B1(new_n253_), .B2(new_n265_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G78gat), .B(G106gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT91), .ZN(new_n349_));
  XOR2_X1   g148(.A(KEYINPUT87), .B(G228gat), .Z(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(G233gat), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT91), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n348_), .B(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(G233gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n347_), .A2(new_n351_), .A3(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n339_), .A2(new_n342_), .A3(new_n316_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n355_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n344_), .A2(new_n356_), .A3(new_n357_), .A4(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n357_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n359_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n358_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n363_));
  OAI22_X1  g162(.A1(new_n361_), .A2(new_n343_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n314_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G15gat), .B(G43gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n232_), .A2(new_n241_), .A3(KEYINPUT30), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT30), .B1(new_n232_), .B2(new_n241_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT30), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n242_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n292_), .A2(KEYINPUT30), .ZN(new_n375_));
  INV_X1    g174(.A(new_n369_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(G71gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(G99gat), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n372_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n372_), .B2(new_n377_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT84), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n381_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n376_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n370_), .A2(new_n371_), .A3(new_n369_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n372_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G134gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G127gat), .ZN(new_n393_));
  INV_X1    g192(.A(G127gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G134gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G113gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(G120gat), .ZN(new_n398_));
  INV_X1    g197(.A(G120gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(G113gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n396_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT31), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n384_), .A2(new_n391_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n388_), .A2(new_n390_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n405_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n384_), .A2(new_n391_), .A3(new_n407_), .A4(new_n405_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G225gat), .A2(G233gat), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n404_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT94), .B(KEYINPUT4), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n396_), .B(new_n402_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n327_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n320_), .A2(new_n322_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n317_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n334_), .A2(new_n328_), .A3(new_n336_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT1), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n318_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n418_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n333_), .A2(new_n337_), .A3(new_n404_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(KEYINPUT4), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n417_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n414_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G1gat), .B(G29gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(G85gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT0), .B(G57gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n434_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n428_), .A2(new_n436_), .A3(new_n429_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n366_), .A2(new_n413_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n365_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n414_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n425_), .A2(new_n426_), .A3(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n442_), .A2(new_n434_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n444_), .A2(KEYINPUT96), .A3(new_n427_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT96), .B1(new_n444_), .B2(new_n427_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n443_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT97), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT97), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n449_), .B(new_n443_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n312_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n437_), .B1(KEYINPUT95), .B2(KEYINPUT33), .ZN(new_n453_));
  NOR2_X1   g252(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n428_), .A2(new_n436_), .A3(new_n429_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n451_), .A2(new_n308_), .A3(new_n452_), .A4(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n305_), .A2(KEYINPUT32), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n295_), .A2(new_n459_), .B1(new_n437_), .B2(new_n435_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n304_), .A2(new_n307_), .A3(new_n458_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n440_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n365_), .A2(new_n438_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n309_), .A2(new_n464_), .A3(new_n313_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n413_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT99), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n413_), .B(KEYINPUT99), .C1(new_n463_), .C2(new_n465_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n439_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G29gat), .B(G36gat), .Z(new_n471_));
  XOR2_X1   g270(.A(G43gat), .B(G50gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475_));
  INV_X1    g274(.A(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G8gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n474_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G229gat), .A2(G233gat), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n473_), .B(KEYINPUT15), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n481_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n474_), .B(new_n481_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n483_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n484_), .A2(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G113gat), .B(G141gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT78), .ZN(new_n491_));
  XOR2_X1   g290(.A(G169gat), .B(G197gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n489_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n470_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G230gat), .A2(G233gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT6), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT64), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT10), .B(G99gat), .Z(new_n506_));
  INV_X1    g305(.A(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G85gat), .B(G92gat), .ZN(new_n510_));
  MUX2_X1   g309(.A(new_n509_), .B(new_n510_), .S(KEYINPUT9), .Z(new_n511_));
  NAND3_X1  g310(.A1(new_n505_), .A2(new_n508_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n510_), .B(KEYINPUT66), .ZN(new_n513_));
  NOR2_X1   g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  AOI211_X1 g315(.A(KEYINPUT8), .B(new_n513_), .C1(new_n505_), .C2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT8), .ZN(new_n518_));
  INV_X1    g317(.A(new_n513_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n500_), .A2(new_n502_), .A3(KEYINPUT67), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n503_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n516_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n518_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n512_), .B1(new_n517_), .B2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G57gat), .B(G64gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT11), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT68), .ZN(new_n528_));
  XOR2_X1   g327(.A(G71gat), .B(G78gat), .Z(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(KEYINPUT11), .B2(new_n526_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n528_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n525_), .A2(new_n532_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n531_), .B(new_n512_), .C1(new_n524_), .C2(new_n517_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(KEYINPUT12), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n525_), .A2(new_n532_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n498_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n497_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G120gat), .B(G148gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G176gat), .B(G204gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(KEYINPUT70), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT13), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT13), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT74), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n531_), .B(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n481_), .B(KEYINPUT73), .Z(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT76), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G127gat), .B(G155gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(G183gat), .B(G211gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n564_), .A2(new_n565_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n558_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT77), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n558_), .A2(new_n566_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n568_), .A2(KEYINPUT77), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n525_), .A2(new_n485_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT34), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT35), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n473_), .B(new_n512_), .C1(new_n517_), .C2(new_n524_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n574_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n577_), .A2(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n574_), .A2(new_n584_), .A3(new_n579_), .A4(new_n580_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT36), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT72), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n589_), .A2(KEYINPUT36), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n583_), .A2(new_n585_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n590_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT72), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n593_), .A2(new_n594_), .A3(new_n597_), .A4(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT37), .B1(new_n596_), .B2(new_n599_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT71), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT71), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n604_), .B(KEYINPUT37), .C1(new_n596_), .C2(new_n599_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n573_), .A2(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n496_), .A2(new_n553_), .A3(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n438_), .B(KEYINPUT100), .Z(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n609_), .A2(new_n476_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n551_), .A2(new_n552_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n615_), .A2(new_n573_), .A3(new_n495_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n593_), .A2(new_n597_), .A3(new_n600_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n470_), .A2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n438_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n612_), .A2(new_n613_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n614_), .A2(new_n623_), .A3(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(new_n314_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n477_), .B1(new_n620_), .B2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT39), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n609_), .A2(new_n477_), .A3(new_n626_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g430(.A(G15gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n413_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n620_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT41), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n609_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1326gat));
  INV_X1    g436(.A(G22gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n365_), .B(KEYINPUT101), .Z(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n609_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n638_), .B1(new_n620_), .B2(new_n640_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT103), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n643_), .A2(new_n644_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n641_), .B1(new_n645_), .B2(new_n646_), .ZN(G1327gat));
  NOR2_X1   g446(.A1(new_n571_), .A2(new_n572_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n615_), .A2(new_n648_), .A3(new_n617_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n496_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n438_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n553_), .A2(new_n494_), .A3(new_n573_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n601_), .A2(new_n603_), .A3(KEYINPUT104), .A4(new_n605_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT43), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n470_), .A2(new_n655_), .A3(new_n606_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(KEYINPUT43), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n633_), .A2(new_n622_), .A3(new_n365_), .A4(new_n314_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n469_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n309_), .A2(new_n464_), .A3(new_n313_), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n448_), .A2(new_n450_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n311_), .A2(new_n312_), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n661_), .A2(new_n662_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n660_), .B1(new_n663_), .B2(new_n440_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT99), .B1(new_n664_), .B2(new_n413_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n658_), .B1(new_n659_), .B2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n657_), .B1(new_n666_), .B2(new_n607_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n653_), .B1(new_n656_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT44), .B1(new_n668_), .B2(KEYINPUT105), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n655_), .B1(new_n470_), .B2(new_n606_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n666_), .A2(new_n607_), .A3(new_n657_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n652_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AOI22_X1  g473(.A1(new_n669_), .A2(new_n674_), .B1(KEYINPUT44), .B2(new_n672_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n611_), .A2(G29gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n651_), .B1(new_n675_), .B2(new_n676_), .ZN(G1328gat));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(KEYINPUT108), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT108), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT109), .Z(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n650_), .A2(new_n683_), .A3(new_n626_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n314_), .B1(new_n672_), .B2(KEYINPUT44), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n688_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT105), .B(new_n652_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G36gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n686_), .B1(new_n692_), .B2(KEYINPUT106), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n691_), .A2(new_n694_), .A3(G36gat), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n679_), .B(new_n682_), .C1(new_n693_), .C2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT44), .B(new_n653_), .C1(new_n656_), .C2(new_n667_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n626_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n669_), .B2(new_n674_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT106), .B1(new_n699_), .B2(new_n683_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n686_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n695_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n679_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n681_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n696_), .A2(new_n704_), .ZN(G1329gat));
  AOI21_X1  g504(.A(G43gat), .B1(new_n650_), .B2(new_n633_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT111), .Z(new_n707_));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n633_), .A2(G43gat), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n675_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n675_), .B2(new_n709_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT47), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n707_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1330gat));
  INV_X1    g515(.A(G50gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n650_), .A2(new_n717_), .A3(new_n640_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n675_), .A2(KEYINPUT112), .A3(new_n440_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G50gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT112), .B1(new_n675_), .B2(new_n440_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(G1331gat));
  NAND4_X1  g521(.A1(new_n619_), .A2(new_n495_), .A3(new_n615_), .A4(new_n648_), .ZN(new_n723_));
  INV_X1    g522(.A(G57gat), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n622_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n470_), .A2(new_n553_), .A3(new_n494_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n608_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n610_), .B1(new_n727_), .B2(KEYINPUT113), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n728_), .B1(KEYINPUT113), .B2(new_n727_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n729_), .B2(new_n724_), .ZN(G1332gat));
  OAI21_X1  g529(.A(G64gat), .B1(new_n723_), .B2(new_n314_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT48), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n314_), .A2(G64gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n727_), .B2(new_n733_), .ZN(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n723_), .B2(new_n413_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT49), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n633_), .A2(new_n379_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n727_), .B2(new_n737_), .ZN(G1334gat));
  OAI21_X1  g537(.A(G78gat), .B1(new_n723_), .B2(new_n639_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT50), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n639_), .A2(G78gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(new_n727_), .B2(new_n741_), .ZN(G1335gat));
  AND3_X1   g541(.A1(new_n726_), .A2(new_n573_), .A3(new_n618_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n611_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT114), .Z(new_n745_));
  NAND2_X1  g544(.A1(new_n670_), .A2(new_n671_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT115), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n615_), .A2(new_n573_), .A3(new_n495_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n438_), .A2(G85gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n745_), .B1(new_n750_), .B2(new_n751_), .ZN(G1336gat));
  OAI21_X1  g551(.A(G92gat), .B1(new_n749_), .B2(new_n314_), .ZN(new_n753_));
  INV_X1    g552(.A(G92gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n743_), .A2(new_n754_), .A3(new_n626_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n749_), .B2(new_n413_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n743_), .A2(new_n633_), .A3(new_n506_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g559(.A1(new_n743_), .A2(new_n507_), .A3(new_n440_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n748_), .A2(new_n365_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n746_), .A2(KEYINPUT116), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G106gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT116), .B1(new_n746_), .B2(new_n762_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n764_), .A2(KEYINPUT52), .A3(new_n765_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n761_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g570(.A1(new_n608_), .A2(new_n495_), .A3(new_n553_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n535_), .A2(new_n537_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n497_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n535_), .A2(new_n498_), .A3(new_n537_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(KEYINPUT55), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n547_), .B1(new_n538_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n489_), .A2(new_n493_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n486_), .A2(new_n482_), .A3(new_n488_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n493_), .B1(new_n487_), .B2(new_n483_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n540_), .B2(new_n545_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n782_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n779_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n789_), .A2(KEYINPUT58), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT120), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT120), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n789_), .A2(new_n794_), .A3(KEYINPUT58), .A4(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n782_), .A2(new_n788_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n790_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n607_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n797_), .B1(new_n607_), .B2(new_n800_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n796_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT121), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n550_), .A2(new_n787_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n546_), .A2(new_n494_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n778_), .A2(new_n781_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT117), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n806_), .B1(new_n808_), .B2(new_n779_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n805_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT118), .B1(new_n811_), .B2(new_n618_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT118), .B(KEYINPUT57), .C1(new_n811_), .C2(new_n618_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n796_), .B(new_n817_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n804_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n774_), .B1(new_n819_), .B2(new_n573_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n366_), .A2(new_n413_), .A3(new_n610_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT59), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n648_), .B1(new_n816_), .B2(new_n803_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n824_), .B(new_n821_), .C1(new_n825_), .C2(new_n774_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n495_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n819_), .A2(new_n573_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n774_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n822_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n397_), .A3(new_n494_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n832_), .ZN(G1340gat));
  OAI211_X1 g632(.A(new_n615_), .B(new_n826_), .C1(new_n831_), .C2(new_n824_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n823_), .A2(KEYINPUT122), .A3(new_n615_), .A4(new_n826_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(G120gat), .A3(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n399_), .B1(new_n553_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n831_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n399_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1341gat));
  OAI21_X1  g640(.A(G127gat), .B1(new_n827_), .B2(new_n573_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n831_), .A2(new_n394_), .A3(new_n648_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1342gat));
  XOR2_X1   g643(.A(KEYINPUT123), .B(G134gat), .Z(new_n845_));
  NOR2_X1   g644(.A1(new_n606_), .A2(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n823_), .A2(new_n826_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G134gat), .B1(new_n831_), .B2(new_n618_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT124), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n848_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  INV_X1    g650(.A(new_n846_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n850_), .B(new_n851_), .C1(new_n827_), .C2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(G1343gat));
  NAND2_X1  g653(.A1(new_n829_), .A2(new_n830_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n626_), .A2(new_n610_), .A3(new_n365_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n413_), .A3(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n495_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n325_), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n553_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n326_), .ZN(G1345gat));
  NOR2_X1   g660(.A1(new_n857_), .A2(new_n573_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT61), .B(G155gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  OAI21_X1  g663(.A(G162gat), .B1(new_n857_), .B2(new_n606_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n617_), .A2(G162gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n857_), .B2(new_n866_), .ZN(G1347gat));
  XNOR2_X1  g666(.A(KEYINPUT22), .B(G169gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n825_), .A2(new_n774_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n611_), .A2(new_n314_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n633_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n639_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n869_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT125), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(KEYINPUT125), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n494_), .B(new_n868_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n878_));
  AOI211_X1 g677(.A(KEYINPUT62), .B(new_n203_), .C1(new_n874_), .C2(new_n494_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n874_), .A2(new_n494_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(G169gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n879_), .B2(new_n882_), .ZN(G1348gat));
  OAI21_X1  g682(.A(new_n615_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n820_), .A2(new_n440_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n553_), .A2(new_n204_), .A3(new_n871_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n884_), .A2(new_n204_), .B1(new_n885_), .B2(new_n886_), .ZN(G1349gat));
  OR2_X1    g686(.A1(new_n869_), .A2(new_n873_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT125), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n875_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n648_), .A2(new_n218_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n885_), .A2(new_n648_), .A3(new_n872_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n891_), .A2(new_n892_), .B1(new_n893_), .B2(new_n214_), .ZN(G1350gat));
  NOR2_X1   g693(.A1(new_n617_), .A2(new_n278_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n891_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n606_), .B1(new_n890_), .B2(new_n875_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n220_), .B2(new_n897_), .ZN(G1351gat));
  AND3_X1   g697(.A1(new_n626_), .A2(new_n413_), .A3(new_n464_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n855_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n495_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n245_), .ZN(G1352gat));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n553_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n248_), .ZN(G1353gat));
  NOR2_X1   g703(.A1(new_n900_), .A2(new_n573_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT63), .B(G211gat), .Z(new_n906_));
  AOI21_X1  g705(.A(KEYINPUT126), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n855_), .A2(new_n648_), .A3(new_n899_), .A4(new_n906_), .ZN(new_n908_));
  OR2_X1    g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n905_), .B2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n907_), .B1(KEYINPUT126), .B2(new_n910_), .ZN(G1354gat));
  XNOR2_X1  g710(.A(KEYINPUT127), .B(G218gat), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n900_), .A2(new_n606_), .A3(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n855_), .A2(new_n618_), .A3(new_n899_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n912_), .ZN(G1355gat));
endmodule


