//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT80), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(KEYINPUT23), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(KEYINPUT23), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(new_n204_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n203_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n213_), .A2(new_n207_), .A3(new_n217_), .A4(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n210_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT30), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G227gat), .A2(G233gat), .ZN(new_n223_));
  INV_X1    g022(.A(G15gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(G43gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G71gat), .B(G99gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n222_), .A2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n229_), .B(KEYINPUT81), .Z(new_n230_));
  NAND2_X1  g029(.A1(new_n222_), .A2(new_n228_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT82), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT84), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n237_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT31), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n233_), .B1(new_n234_), .B2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n234_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n213_), .A2(new_n219_), .A3(new_n217_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n208_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT91), .ZN(new_n249_));
  XOR2_X1   g048(.A(G197gat), .B(G204gat), .Z(new_n250_));
  OR2_X1    g049(.A1(new_n250_), .A2(KEYINPUT21), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(KEYINPUT21), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n252_), .A2(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n207_), .B1(G183gat), .B2(G190gat), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n257_), .A2(new_n203_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n249_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n221_), .A2(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G226gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT19), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT20), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n260_), .A2(new_n261_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT92), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT92), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n260_), .A2(new_n268_), .A3(new_n261_), .A4(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT91), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n248_), .B(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n256_), .B1(new_n272_), .B2(new_n258_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n221_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n256_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n264_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n263_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT18), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G64gat), .B(G92gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n270_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n256_), .A2(new_n258_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT20), .B1(new_n284_), .B2(new_n248_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n261_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n263_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(new_n277_), .B2(new_n263_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n282_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n283_), .A2(new_n290_), .A3(KEYINPUT27), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n283_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n282_), .B1(new_n270_), .B2(new_n278_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT27), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n292_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n299_), .B1(new_n302_), .B2(KEYINPUT1), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(KEYINPUT1), .B2(new_n302_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n306_), .B(KEYINPUT3), .Z(new_n309_));
  XOR2_X1   g108(.A(new_n305_), .B(KEYINPUT2), .Z(new_n310_));
  OAI221_X1 g109(.A(new_n302_), .B1(G155gat), .B2(G162gat), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n240_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT93), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n308_), .A2(new_n239_), .A3(new_n238_), .A4(new_n311_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  OR3_X1    g115(.A1(new_n312_), .A2(new_n314_), .A3(new_n240_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT4), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G225gat), .A2(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n312_), .A2(new_n322_), .A3(new_n240_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT94), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n319_), .A2(new_n321_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT96), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G1gat), .B(G29gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT95), .B(G85gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT0), .B(G57gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n318_), .A2(new_n327_), .A3(new_n320_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n326_), .A2(new_n329_), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI211_X1 g137(.A(KEYINPUT96), .B(new_n321_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n328_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n335_), .B1(new_n340_), .B2(new_n326_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G22gat), .B(G50gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n312_), .A2(KEYINPUT29), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT28), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n312_), .A2(KEYINPUT29), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n344_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n346_), .A2(new_n349_), .A3(new_n344_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n353_), .A2(KEYINPUT90), .ZN(new_n356_));
  INV_X1    g155(.A(new_n349_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n347_), .A2(new_n348_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n357_), .A2(new_n358_), .A3(new_n343_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n356_), .B1(new_n359_), .B2(new_n350_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(KEYINPUT88), .A2(KEYINPUT29), .ZN(new_n362_));
  AND2_X1   g161(.A1(KEYINPUT88), .A2(KEYINPUT29), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n312_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n275_), .B1(new_n364_), .B2(KEYINPUT89), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(KEYINPUT89), .B2(new_n364_), .ZN(new_n366_));
  INV_X1    g165(.A(G228gat), .ZN(new_n367_));
  OR2_X1    g166(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  AOI211_X1 g170(.A(new_n275_), .B(new_n370_), .C1(new_n312_), .C2(KEYINPUT29), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT87), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n361_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n355_), .A2(new_n374_), .A3(new_n360_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n298_), .A2(new_n342_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT97), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(KEYINPUT33), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n337_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n340_), .A2(new_n335_), .A3(new_n326_), .A4(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n318_), .A2(KEYINPUT98), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n318_), .A2(KEYINPUT98), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n321_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n319_), .A2(new_n320_), .A3(new_n325_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n334_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n382_), .A2(new_n295_), .A3(new_n384_), .A4(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n288_), .A2(KEYINPUT32), .A3(new_n282_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n270_), .A2(new_n278_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n282_), .A2(KEYINPUT32), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n378_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n379_), .B1(new_n396_), .B2(KEYINPUT99), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT99), .ZN(new_n398_));
  AOI211_X1 g197(.A(new_n398_), .B(new_n378_), .C1(new_n390_), .C2(new_n395_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n246_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n298_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n401_), .A2(new_n246_), .A3(new_n378_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n342_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G29gat), .B(G36gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT70), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G43gat), .B(G50gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT70), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n405_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT15), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n408_), .A2(new_n412_), .A3(KEYINPUT15), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT73), .B(G15gat), .ZN(new_n418_));
  INV_X1    g217(.A(G22gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G1gat), .ZN(new_n421_));
  INV_X1    g220(.A(G8gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT14), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(G1gat), .B(G8gat), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n420_), .A2(new_n425_), .A3(new_n423_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n417_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G229gat), .A2(G233gat), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n427_), .A2(new_n408_), .A3(new_n412_), .A4(new_n428_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n428_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n425_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n413_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT78), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n429_), .A2(KEYINPUT78), .A3(new_n413_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n433_), .B1(new_n440_), .B2(new_n431_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G113gat), .B(G141gat), .Z(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT79), .ZN(new_n443_));
  XOR2_X1   g242(.A(G169gat), .B(G197gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n445_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n404_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G230gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  OR2_X1    g250(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n452_));
  INV_X1    g251(.A(G106gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT64), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n462_), .B1(new_n456_), .B2(new_n455_), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G85gat), .A2(G92gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(KEYINPUT9), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT9), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(G85gat), .A3(G92gat), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n457_), .B(new_n463_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT8), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n458_), .A2(KEYINPUT68), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT68), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n480_));
  NOR2_X1   g279(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n476_), .B(new_n478_), .C1(new_n481_), .C2(new_n480_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(G99gat), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n487_), .B(new_n453_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(new_n484_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n466_), .A2(new_n467_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n475_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n462_), .ZN(new_n494_));
  AOI211_X1 g293(.A(KEYINPUT8), .B(new_n491_), .C1(new_n494_), .C2(new_n489_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n474_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n498_));
  XOR2_X1   g297(.A(G71gat), .B(G78gat), .Z(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n499_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n496_), .A2(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n474_), .B(new_n503_), .C1(new_n493_), .C2(new_n495_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(KEYINPUT12), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(KEYINPUT12), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n494_), .A2(new_n489_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n475_), .A3(new_n492_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n479_), .A2(new_n482_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n491_), .B1(new_n511_), .B2(new_n484_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n512_), .B2(new_n475_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n503_), .B1(new_n513_), .B2(new_n474_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n508_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n451_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n450_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G120gat), .B(G148gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT5), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G176gat), .B(G204gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n522_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(KEYINPUT69), .B(new_n522_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT13), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n429_), .B(KEYINPUT74), .Z(new_n533_));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT75), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n503_), .B(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n536_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G127gat), .B(G155gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G183gat), .B(G211gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT17), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n544_), .B(KEYINPUT17), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n537_), .A2(new_n547_), .A3(new_n538_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT77), .Z(new_n550_));
  AOI22_X1  g349(.A1(new_n415_), .A2(new_n416_), .B1(new_n513_), .B2(new_n474_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G232gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT34), .ZN(new_n553_));
  OAI22_X1  g352(.A1(new_n496_), .A2(new_n413_), .B1(KEYINPUT35), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT35), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OR3_X1    g356(.A1(new_n551_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n551_), .B2(new_n554_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(KEYINPUT72), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT71), .ZN(new_n562_));
  XOR2_X1   g361(.A(G134gat), .B(G162gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n560_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n558_), .A2(KEYINPUT72), .A3(new_n559_), .A4(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n558_), .A2(new_n559_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT36), .A3(new_n564_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT37), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT37), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n569_), .A2(new_n574_), .A3(new_n571_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n550_), .A2(new_n576_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n449_), .A2(new_n532_), .A3(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n342_), .A2(KEYINPUT100), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n342_), .A2(KEYINPUT100), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(new_n421_), .A3(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT38), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n572_), .B(KEYINPUT101), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT102), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n531_), .A2(new_n549_), .A3(new_n448_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT103), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n342_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n583_), .B1(new_n421_), .B2(new_n594_), .ZN(G1324gat));
  NAND3_X1  g394(.A1(new_n578_), .A2(new_n422_), .A3(new_n401_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT104), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n587_), .A2(new_n598_), .A3(new_n401_), .A4(new_n589_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(G8gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n587_), .A2(new_n401_), .A3(new_n589_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT104), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n597_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  AND4_X1   g402(.A1(new_n597_), .A2(new_n602_), .A3(G8gat), .A4(new_n599_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n596_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(G1325gat));
  NAND3_X1  g406(.A1(new_n578_), .A2(new_n224_), .A3(new_n245_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n592_), .A2(new_n245_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n609_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT41), .B1(new_n609_), .B2(G15gat), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n608_), .B1(new_n610_), .B2(new_n611_), .ZN(G1326gat));
  XNOR2_X1  g411(.A(new_n378_), .B(KEYINPUT105), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n578_), .A2(new_n419_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n592_), .A2(new_n614_), .ZN(new_n616_));
  XOR2_X1   g415(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n617_));
  AND3_X1   g416(.A1(new_n616_), .A2(G22gat), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n616_), .B2(G22gat), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(G1327gat));
  INV_X1    g419(.A(new_n448_), .ZN(new_n621_));
  OR3_X1    g420(.A1(new_n532_), .A2(new_n621_), .A3(new_n550_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT43), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n573_), .A2(new_n575_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n404_), .B2(new_n625_), .ZN(new_n626_));
  AOI211_X1 g425(.A(KEYINPUT43), .B(new_n576_), .C1(new_n400_), .C2(new_n403_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT44), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI211_X1 g429(.A(KEYINPUT44), .B(new_n623_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n630_), .A2(G29gat), .A3(new_n581_), .A4(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(G29gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n584_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n634_), .A2(new_n532_), .A3(new_n550_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n404_), .A2(new_n448_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT107), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n404_), .A2(new_n638_), .A3(new_n448_), .A4(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n633_), .B1(new_n640_), .B2(new_n342_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n632_), .A2(new_n641_), .ZN(G1328gat));
  NAND3_X1  g441(.A1(new_n630_), .A2(new_n401_), .A3(new_n631_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G36gat), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n298_), .A2(G36gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n637_), .A2(new_n639_), .A3(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT45), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT46), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n644_), .A2(KEYINPUT46), .A3(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1329gat));
  NAND4_X1  g451(.A1(new_n630_), .A2(G43gat), .A3(new_n245_), .A4(new_n631_), .ZN(new_n653_));
  INV_X1    g452(.A(G43gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n654_), .B1(new_n640_), .B2(new_n246_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g456(.A1(new_n630_), .A2(G50gat), .A3(new_n378_), .A4(new_n631_), .ZN(new_n658_));
  INV_X1    g457(.A(G50gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n659_), .B1(new_n640_), .B2(new_n613_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n658_), .A2(new_n660_), .ZN(G1331gat));
  NOR2_X1   g460(.A1(new_n531_), .A2(new_n448_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n587_), .A2(new_n550_), .A3(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(KEYINPUT109), .A2(G57gat), .ZN(new_n664_));
  AND2_X1   g463(.A1(KEYINPUT109), .A2(G57gat), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n663_), .B(new_n593_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n404_), .A2(new_n621_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT108), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n531_), .B1(new_n667_), .B2(KEYINPUT108), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n581_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n670_), .A2(new_n577_), .A3(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n666_), .B1(new_n672_), .B2(G57gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT110), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT110), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n675_), .B(new_n666_), .C1(new_n672_), .C2(G57gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1332gat));
  INV_X1    g476(.A(G64gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n663_), .B2(new_n401_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT48), .Z(new_n680_));
  OR2_X1    g479(.A1(new_n670_), .A2(new_n577_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n401_), .A2(new_n678_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n680_), .B1(new_n681_), .B2(new_n682_), .ZN(G1333gat));
  INV_X1    g482(.A(G71gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n663_), .B2(new_n245_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT49), .Z(new_n686_));
  NAND2_X1  g485(.A1(new_n245_), .A2(new_n684_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n681_), .B2(new_n687_), .ZN(G1334gat));
  NAND2_X1  g487(.A1(new_n663_), .A2(new_n614_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G78gat), .ZN(new_n690_));
  XOR2_X1   g489(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n613_), .A2(G78gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n681_), .B2(new_n693_), .ZN(G1335gat));
  NOR3_X1   g493(.A1(new_n550_), .A2(new_n531_), .A3(new_n448_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G85gat), .B1(new_n696_), .B2(new_n342_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n634_), .A2(new_n550_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n668_), .A2(new_n698_), .A3(new_n669_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n581_), .A2(new_n464_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(G1336gat));
  OAI21_X1  g500(.A(G92gat), .B1(new_n696_), .B2(new_n298_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n401_), .A2(new_n465_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n699_), .B2(new_n703_), .ZN(G1337gat));
  OAI21_X1  g503(.A(G99gat), .B1(new_n696_), .B2(new_n246_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n245_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n699_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g507(.A(new_n378_), .B(new_n695_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710_));
  AND4_X1   g509(.A1(KEYINPUT112), .A2(new_n709_), .A3(new_n710_), .A4(G106gat), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n453_), .B1(new_n712_), .B2(KEYINPUT52), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n709_), .A2(new_n713_), .B1(KEYINPUT112), .B2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n378_), .A2(new_n453_), .ZN(new_n715_));
  OAI22_X1  g514(.A1(new_n711_), .A2(new_n714_), .B1(new_n699_), .B2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  OAI221_X1 g518(.A(new_n717_), .B1(new_n699_), .B2(new_n715_), .C1(new_n711_), .C2(new_n714_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1339gat));
  NAND4_X1  g520(.A1(new_n576_), .A2(new_n550_), .A3(new_n531_), .A4(new_n621_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT54), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT116), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n508_), .A2(new_n514_), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT12), .B(new_n503_), .C1(new_n513_), .C2(new_n474_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT55), .B(new_n450_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n507_), .A2(new_n515_), .A3(new_n451_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n507_), .A2(new_n515_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT55), .B1(new_n732_), .B2(new_n450_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n522_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT56), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT114), .B(new_n522_), .C1(new_n731_), .C2(new_n733_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n736_), .A2(KEYINPUT115), .A3(new_n737_), .A4(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n448_), .A2(new_n524_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT56), .B(new_n522_), .C1(new_n731_), .C2(new_n733_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT56), .B1(new_n734_), .B2(new_n735_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n738_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n726_), .B1(new_n741_), .B2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n744_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n750_), .A2(KEYINPUT116), .A3(new_n739_), .A4(new_n740_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n438_), .A2(new_n431_), .A3(new_n439_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n445_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(KEYINPUT117), .A3(new_n445_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n430_), .A2(G229gat), .A3(G233gat), .A4(new_n432_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n446_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(new_n528_), .A3(new_n527_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n747_), .A2(new_n751_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT57), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n584_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n734_), .A2(new_n737_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n742_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n446_), .A2(new_n758_), .A3(new_n524_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(KEYINPUT58), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n625_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT58), .B1(new_n766_), .B2(new_n767_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n764_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT57), .B1(new_n761_), .B2(new_n634_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n725_), .B1(new_n775_), .B2(new_n550_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n402_), .A2(new_n581_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT59), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n549_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n725_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n777_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n784_), .B2(new_n778_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n777_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n788_), .A2(KEYINPUT59), .B1(new_n776_), .B2(new_n779_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT118), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n448_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G113gat), .ZN(new_n792_));
  OR3_X1    g591(.A1(new_n788_), .A2(G113gat), .A3(new_n621_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1340gat));
  INV_X1    g593(.A(G120gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n531_), .B2(KEYINPUT60), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n784_), .B(new_n796_), .C1(KEYINPUT60), .C2(new_n795_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n789_), .A2(new_n532_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n797_), .B1(new_n799_), .B2(new_n795_), .ZN(G1341gat));
  INV_X1    g599(.A(G127gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n784_), .A2(new_n801_), .A3(new_n550_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n787_), .A2(new_n549_), .A3(new_n790_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n801_), .ZN(G1342gat));
  NAND3_X1  g603(.A1(new_n787_), .A2(new_n625_), .A3(new_n790_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(G134gat), .ZN(new_n806_));
  OR3_X1    g605(.A1(new_n788_), .A2(G134gat), .A3(new_n585_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1343gat));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  INV_X1    g608(.A(new_n378_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n245_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n782_), .B2(new_n725_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n581_), .A2(new_n298_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n809_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n771_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n760_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n750_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n726_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n584_), .B1(new_n820_), .B2(new_n751_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n817_), .B1(new_n821_), .B2(KEYINPUT57), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n724_), .B1(new_n822_), .B2(new_n781_), .ZN(new_n823_));
  NOR4_X1   g622(.A1(new_n823_), .A2(KEYINPUT119), .A3(new_n812_), .A4(new_n814_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n448_), .B1(new_n816_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT121), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n761_), .A2(new_n634_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n762_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n549_), .B1(new_n828_), .B2(new_n817_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n811_), .B(new_n815_), .C1(new_n829_), .C2(new_n724_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT119), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n783_), .A2(new_n809_), .A3(new_n811_), .A4(new_n815_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n448_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT120), .B(G141gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n826_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n836_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n834_), .B1(new_n833_), .B2(new_n448_), .ZN(new_n839_));
  AOI211_X1 g638(.A(KEYINPUT121), .B(new_n621_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n837_), .A2(new_n841_), .ZN(G1344gat));
  NAND2_X1  g641(.A1(new_n833_), .A2(new_n532_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g643(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT61), .B(G155gat), .Z(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n833_), .A2(new_n550_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n833_), .B2(new_n550_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n846_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n851_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n845_), .A3(new_n849_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1346gat));
  INV_X1    g654(.A(new_n833_), .ZN(new_n856_));
  OR3_X1    g655(.A1(new_n856_), .A2(G162gat), .A3(new_n585_), .ZN(new_n857_));
  OAI21_X1  g656(.A(G162gat), .B1(new_n856_), .B2(new_n576_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1347gat));
  NOR2_X1   g658(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n401_), .A2(new_n245_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n614_), .A2(new_n581_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n776_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n621_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n214_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n860_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NOR4_X1   g666(.A1(new_n864_), .A2(KEYINPUT124), .A3(KEYINPUT62), .A4(new_n214_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT22), .B(G169gat), .Z(new_n869_));
  OAI22_X1  g668(.A1(new_n867_), .A2(new_n868_), .B1(new_n865_), .B2(new_n869_), .ZN(G1348gat));
  INV_X1    g669(.A(new_n863_), .ZN(new_n871_));
  AOI21_X1  g670(.A(G176gat), .B1(new_n871_), .B2(new_n532_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n823_), .A2(new_n378_), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n581_), .A2(new_n861_), .A3(new_n215_), .A4(new_n531_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(G1349gat));
  OR3_X1    g674(.A1(new_n863_), .A2(new_n211_), .A3(new_n781_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n877_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n581_), .A2(new_n861_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n880_), .A2(new_n550_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G183gat), .B1(new_n873_), .B2(new_n881_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n878_), .A2(new_n879_), .A3(new_n882_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n863_), .B2(new_n576_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n586_), .A2(new_n212_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n863_), .B2(new_n885_), .ZN(G1351gat));
  NAND3_X1  g685(.A1(new_n813_), .A2(new_n342_), .A3(new_n401_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n621_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n531_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT126), .B(G204gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1353gat));
  NOR2_X1   g691(.A1(new_n887_), .A2(new_n781_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n893_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT63), .B(G211gat), .Z(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n893_), .B2(new_n895_), .ZN(G1354gat));
  INV_X1    g695(.A(G218gat), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n887_), .A2(new_n897_), .A3(new_n576_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n887_), .A2(KEYINPUT127), .A3(new_n585_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(G218gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT127), .B1(new_n887_), .B2(new_n585_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n898_), .B1(new_n900_), .B2(new_n901_), .ZN(G1355gat));
endmodule


