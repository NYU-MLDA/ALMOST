//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G78gat), .Z(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n204_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT7), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  INV_X1    g022(.A(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n221_), .A2(new_n222_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n217_), .A2(KEYINPUT66), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT6), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n216_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n213_), .A2(new_n214_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n232_), .A3(new_n216_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n227_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n229_), .B1(new_n237_), .B2(new_n222_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239_));
  OR2_X1    g038(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n212_), .A3(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n225_), .A2(KEYINPUT9), .A3(new_n226_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT9), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(G85gat), .A3(G92gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n218_), .A2(new_n246_), .A3(new_n219_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n239_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n247_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n249_), .A2(KEYINPUT65), .A3(new_n242_), .A4(new_n243_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n209_), .B1(new_n238_), .B2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n230_), .A2(new_n232_), .A3(new_n216_), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n253_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT8), .B1(new_n254_), .B2(new_n227_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n255_), .A2(new_n229_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n209_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n257_), .B2(KEYINPUT67), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(KEYINPUT67), .B2(new_n257_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT64), .Z(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n252_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n252_), .A2(KEYINPUT12), .ZN(new_n267_));
  INV_X1    g066(.A(new_n265_), .ZN(new_n268_));
  OAI211_X1 g067(.A(KEYINPUT69), .B(new_n268_), .C1(new_n256_), .C2(new_n209_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n262_), .B1(new_n256_), .B2(new_n209_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n230_), .A2(new_n232_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n216_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(new_n215_), .A3(new_n236_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n222_), .B1(new_n277_), .B2(new_n228_), .ZN(new_n278_));
  AOI211_X1 g077(.A(KEYINPUT8), .B(new_n227_), .C1(new_n215_), .C2(new_n220_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n251_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n207_), .A2(new_n208_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(new_n205_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n265_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n283_), .A2(KEYINPUT69), .B1(new_n252_), .B2(KEYINPUT12), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n284_), .A2(KEYINPUT70), .A3(new_n266_), .A4(new_n270_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G120gat), .B(G148gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT5), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G176gat), .B(G204gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n263_), .A2(new_n273_), .A3(new_n285_), .A4(new_n289_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n263_), .A2(new_n273_), .A3(new_n285_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n289_), .B(KEYINPUT71), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n296_));
  OAI21_X1  g095(.A(new_n295_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT14), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT77), .B(G8gat), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(G1gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT78), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G15gat), .B(G22gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G231gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n209_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n308_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G127gat), .B(G155gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT16), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G183gat), .B(G211gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT17), .Z(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT81), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n313_), .A2(new_n321_), .A3(new_n318_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(KEYINPUT17), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT79), .Z(new_n324_));
  AOI22_X1  g123(.A1(new_n320_), .A2(new_n322_), .B1(new_n311_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G43gat), .B(G50gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G29gat), .B(G36gat), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(KEYINPUT73), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(KEYINPUT73), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n326_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n328_), .A2(new_n329_), .A3(new_n326_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(new_n238_), .A3(new_n251_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT15), .ZN(new_n335_));
  INV_X1    g134(.A(new_n332_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n335_), .B1(new_n336_), .B2(new_n330_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n331_), .A2(KEYINPUT15), .A3(new_n332_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n334_), .B1(new_n339_), .B2(new_n256_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G232gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT34), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n342_), .A2(KEYINPUT35), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(KEYINPUT35), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(KEYINPUT75), .A3(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n334_), .B(new_n343_), .C1(new_n339_), .C2(new_n256_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT75), .B1(new_n340_), .B2(new_n345_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G190gat), .B(G218gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G134gat), .B(G162gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(KEYINPUT36), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n351_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n340_), .A2(new_n345_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n359_), .A2(new_n351_), .A3(new_n347_), .A4(new_n346_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n355_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n347_), .A3(new_n346_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n354_), .A2(KEYINPUT36), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n356_), .A2(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT37), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n366_), .A2(new_n367_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n363_), .A2(new_n364_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n355_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n360_), .A2(new_n361_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n372_), .B(new_n368_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n369_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n297_), .A2(new_n325_), .A3(new_n371_), .A4(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT103), .ZN(new_n378_));
  XOR2_X1   g177(.A(G211gat), .B(G218gat), .Z(new_n379_));
  INV_X1    g178(.A(G204gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G197gat), .ZN(new_n381_));
  INV_X1    g180(.A(G197gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G204gat), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(KEYINPUT91), .B(KEYINPUT21), .Z(new_n385_));
  AOI21_X1  g184(.A(new_n379_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT90), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n380_), .A3(G197gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n383_), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT21), .B(new_n388_), .C1(new_n389_), .C2(new_n387_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n379_), .A2(KEYINPUT21), .A3(new_n389_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(G233gat), .ZN(new_n394_));
  OR2_X1    g193(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G155gat), .B(G162gat), .Z(new_n399_));
  INV_X1    g198(.A(G141gat), .ZN(new_n400_));
  INV_X1    g199(.A(G148gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT3), .ZN(new_n403_));
  OR3_X1    g202(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G141gat), .A2(G148gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT88), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n403_), .B(new_n404_), .C1(KEYINPUT2), .C2(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n407_), .A2(KEYINPUT2), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n399_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT1), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n399_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n412_), .A2(new_n405_), .A3(new_n402_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT29), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n398_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n398_), .A2(KEYINPUT92), .A3(new_n416_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n391_), .A2(new_n392_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT93), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n416_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n397_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G78gat), .B(G106gat), .Z(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n428_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n421_), .A2(new_n430_), .A3(new_n426_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n415_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT28), .ZN(new_n436_));
  XOR2_X1   g235(.A(G22gat), .B(G50gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n432_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G8gat), .B(G36gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT18), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT32), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G183gat), .A2(G190gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT23), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G169gat), .ZN(new_n453_));
  INV_X1    g252(.A(G176gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n455_), .A2(KEYINPUT24), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT25), .B(G183gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT26), .B(G190gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G169gat), .A2(G176gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n455_), .A2(KEYINPUT24), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(KEYINPUT94), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT94), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n452_), .B(new_n456_), .C1(new_n463_), .C2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT22), .B(G169gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n454_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n450_), .B(new_n451_), .C1(G183gat), .C2(G190gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT95), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n460_), .B(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT96), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n393_), .B1(new_n466_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT19), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT84), .B1(new_n453_), .B2(KEYINPUT22), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT22), .ZN(new_n479_));
  AOI21_X1  g278(.A(G176gat), .B1(new_n479_), .B2(G169gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n453_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n469_), .B(new_n460_), .C1(new_n478_), .C2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n459_), .A2(new_n452_), .A3(new_n456_), .A4(new_n461_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT20), .B1(new_n422_), .B2(new_n485_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n474_), .A2(new_n477_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n466_), .A2(new_n473_), .A3(new_n393_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT20), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n422_), .B2(new_n485_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n476_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n447_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G29gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(G85gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT0), .B(G57gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G127gat), .B(G134gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G113gat), .B(G120gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n415_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n410_), .A2(new_n414_), .A3(new_n500_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(KEYINPUT4), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT4), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n415_), .A2(new_n505_), .A3(new_n501_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n497_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n508_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n514_), .A2(new_n496_), .A3(new_n511_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n492_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n447_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n466_), .A2(new_n472_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n424_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n422_), .B2(new_n485_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n477_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n474_), .A2(new_n476_), .A3(new_n486_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n517_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT102), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT102), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(new_n517_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n516_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n491_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n486_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n466_), .A2(new_n473_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n476_), .B(new_n530_), .C1(new_n531_), .C2(new_n393_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n446_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n446_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT97), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT97), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n529_), .A2(new_n532_), .A3(new_n537_), .A4(new_n533_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n496_), .B1(new_n514_), .B2(new_n511_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT33), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT98), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n540_), .B(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n502_), .A2(new_n509_), .A3(new_n503_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n497_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n545_), .A2(KEYINPUT99), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(KEYINPUT99), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n546_), .B(new_n547_), .C1(new_n509_), .C2(new_n507_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n539_), .A2(new_n543_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n528_), .B1(new_n549_), .B2(KEYINPUT100), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT100), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n539_), .A2(new_n543_), .A3(new_n551_), .A4(new_n548_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n442_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n513_), .A2(new_n515_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n442_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT27), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n536_), .A2(new_n556_), .A3(new_n538_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n533_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT27), .A3(new_n535_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n553_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G227gat), .A2(G233gat), .ZN(new_n563_));
  INV_X1    g362(.A(G15gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(G71gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n483_), .A2(new_n484_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT30), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(G99gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n485_), .B(KEYINPUT30), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n211_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT85), .B(G43gat), .Z(new_n573_));
  AND3_X1   g372(.A1(new_n570_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n567_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n570_), .A2(new_n572_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n573_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n570_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n566_), .A3(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n576_), .A2(new_n581_), .A3(KEYINPUT87), .ZN(new_n582_));
  XOR2_X1   g381(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n583_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n576_), .A2(new_n581_), .A3(KEYINPUT87), .A4(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n501_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n584_), .A2(new_n501_), .A3(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n378_), .B1(new_n562_), .B2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n442_), .A2(new_n560_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n592_), .A3(new_n554_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n584_), .A2(new_n501_), .A3(new_n586_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(new_n587_), .ZN(new_n595_));
  OAI211_X1 g394(.A(KEYINPUT103), .B(new_n595_), .C1(new_n553_), .C2(new_n561_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n591_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n307_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n304_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n336_), .A2(new_n330_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n333_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n599_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n339_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n607_), .A3(new_n598_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G113gat), .B(G141gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G169gat), .B(G197gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n610_), .B(new_n611_), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT82), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n609_), .B(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT83), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT104), .B1(new_n597_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n597_), .A2(KEYINPUT104), .A3(new_n617_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n377_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(G1gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n554_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT38), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n549_), .A2(KEYINPUT100), .ZN(new_n627_));
  INV_X1    g426(.A(new_n528_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(new_n552_), .A3(new_n628_), .ZN(new_n629_));
  OAI22_X1  g428(.A1(new_n629_), .A2(new_n442_), .B1(new_n560_), .B2(new_n555_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT103), .B1(new_n630_), .B2(new_n595_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n596_), .A2(new_n593_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n325_), .B(new_n365_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n615_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n297_), .A2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT105), .Z(new_n636_));
  NOR2_X1   g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n622_), .B1(new_n637_), .B2(new_n623_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n626_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n625_), .B2(new_n624_), .ZN(G1324gat));
  INV_X1    g439(.A(new_n299_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n621_), .A2(new_n560_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n637_), .A2(new_n560_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G8gat), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(KEYINPUT39), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(KEYINPUT39), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n647_), .B(new_n648_), .Z(G1325gat));
  AOI21_X1  g448(.A(new_n564_), .B1(new_n637_), .B2(new_n590_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT41), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n621_), .A2(new_n564_), .A3(new_n590_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1326gat));
  INV_X1    g452(.A(G22gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n637_), .B2(new_n442_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT42), .Z(new_n656_));
  NAND3_X1  g455(.A1(new_n621_), .A2(new_n654_), .A3(new_n442_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1327gat));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(KEYINPUT107), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n376_), .A2(new_n371_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n659_), .A2(KEYINPUT107), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n660_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT43), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n666_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n591_), .A2(new_n665_), .A3(new_n593_), .A4(new_n596_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n661_), .A3(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n664_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n636_), .A2(new_n325_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT44), .A3(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n664_), .A2(new_n669_), .A3(new_n671_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(new_n623_), .A3(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n325_), .A2(new_n365_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n297_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n554_), .A2(G29gat), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n676_), .A2(G29gat), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT109), .ZN(G1328gat));
  NAND3_X1  g481(.A1(new_n672_), .A2(new_n560_), .A3(new_n675_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G36gat), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT110), .ZN(new_n685_));
  AOI21_X1  g484(.A(G36gat), .B1(new_n557_), .B2(new_n559_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n679_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n678_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n620_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n688_), .B(new_n686_), .C1(new_n689_), .C2(new_n618_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT110), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n687_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n687_), .A2(KEYINPUT45), .A3(new_n691_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n684_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n684_), .A2(new_n694_), .A3(KEYINPUT46), .A4(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  AND4_X1   g499(.A1(G43gat), .A2(new_n672_), .A3(new_n590_), .A4(new_n675_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n679_), .A2(new_n590_), .ZN(new_n704_));
  INV_X1    g503(.A(G43gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT111), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n704_), .A2(KEYINPUT111), .A3(new_n705_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n702_), .B(new_n703_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n706_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT47), .B1(new_n709_), .B2(new_n701_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n679_), .B2(new_n442_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n672_), .A2(new_n675_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n442_), .A2(G50gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(G1331gat));
  NOR3_X1   g514(.A1(new_n633_), .A2(new_n617_), .A3(new_n297_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n554_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n597_), .A2(new_n615_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n297_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n325_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(new_n661_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n719_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(G57gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n623_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n718_), .A2(new_n725_), .ZN(G1332gat));
  INV_X1    g525(.A(G64gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n723_), .A2(new_n727_), .A3(new_n560_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n716_), .A2(new_n560_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G64gat), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(KEYINPUT48), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(KEYINPUT48), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT112), .ZN(G1333gat));
  INV_X1    g533(.A(G71gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n716_), .B2(new_n590_), .ZN(new_n736_));
  XOR2_X1   g535(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n723_), .A2(new_n735_), .A3(new_n590_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1334gat));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n716_), .B2(new_n442_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT50), .Z(new_n743_));
  NAND2_X1  g542(.A1(new_n442_), .A2(new_n741_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT114), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n723_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(G1335gat));
  AND3_X1   g546(.A1(new_n719_), .A2(new_n720_), .A3(new_n677_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(new_n223_), .A3(new_n623_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n720_), .A2(new_n721_), .A3(new_n615_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT115), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n670_), .A2(new_n751_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n752_), .A2(KEYINPUT116), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(KEYINPUT116), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(new_n623_), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n749_), .B1(new_n755_), .B2(new_n223_), .ZN(G1336gat));
  NAND3_X1  g555(.A1(new_n748_), .A2(new_n224_), .A3(new_n560_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n753_), .A2(new_n560_), .A3(new_n754_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(new_n224_), .ZN(G1337gat));
  NAND3_X1  g558(.A1(new_n670_), .A2(new_n590_), .A3(new_n751_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n590_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n760_), .A2(G99gat), .B1(new_n748_), .B2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n764_), .B(new_n765_), .ZN(G1338gat));
  NAND4_X1  g565(.A1(new_n664_), .A2(new_n669_), .A3(new_n442_), .A4(new_n751_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G106gat), .B1(new_n767_), .B2(new_n768_), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT52), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n670_), .A2(KEYINPUT118), .A3(new_n442_), .A4(new_n751_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n767_), .A2(new_n768_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n772_), .A2(new_n773_), .A3(G106gat), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n771_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n748_), .A2(new_n212_), .A3(new_n442_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n776_), .A2(new_n780_), .A3(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1339gat));
  AND3_X1   g581(.A1(new_n590_), .A2(new_n592_), .A3(new_n623_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n634_), .A2(new_n290_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n273_), .A2(new_n285_), .A3(new_n785_), .ZN(new_n786_));
  AND4_X1   g585(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .A4(new_n257_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n787_), .A2(KEYINPUT55), .B1(new_n788_), .B2(new_n262_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n292_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n292_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT119), .B1(new_n790_), .B2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n792_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n794_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT119), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n784_), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n598_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n606_), .A2(new_n607_), .A3(new_n599_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n612_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n613_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT120), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n613_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n606_), .A2(new_n607_), .A3(new_n598_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n306_), .A2(new_n333_), .A3(new_n307_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n598_), .B1(new_n607_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n612_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n807_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n293_), .A2(new_n805_), .A3(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT57), .B(new_n365_), .C1(new_n800_), .C2(new_n814_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n813_), .A2(new_n805_), .A3(new_n290_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n792_), .B2(new_n798_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n816_), .B(KEYINPUT58), .C1(new_n792_), .C2(new_n798_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n661_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n815_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n790_), .A2(new_n791_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n793_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n273_), .A2(new_n785_), .A3(new_n285_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n788_), .A2(new_n262_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n785_), .B2(new_n271_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n794_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n824_), .A2(new_n830_), .A3(new_n799_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n784_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n814_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n365_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT121), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n837_), .B(new_n365_), .C1(new_n800_), .C2(new_n814_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n836_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n822_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n835_), .A2(new_n838_), .A3(KEYINPUT122), .A4(new_n836_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n325_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n722_), .A2(new_n844_), .A3(new_n616_), .A4(new_n297_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT54), .B1(new_n377_), .B2(new_n617_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n783_), .B1(new_n843_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n815_), .A2(new_n821_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n839_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n847_), .B1(new_n852_), .B2(new_n721_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n783_), .A2(new_n850_), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n849_), .A2(new_n850_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n616_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n615_), .A2(G113gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n848_), .B2(new_n857_), .ZN(G1340gat));
  NOR2_X1   g657(.A1(new_n297_), .A2(KEYINPUT60), .ZN(new_n859_));
  MUX2_X1   g658(.A(new_n859_), .B(KEYINPUT60), .S(G120gat), .Z(new_n860_));
  NAND2_X1  g659(.A1(new_n849_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n720_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n848_), .B2(KEYINPUT59), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  OAI21_X1  g663(.A(G120gat), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  AOI211_X1 g664(.A(KEYINPUT123), .B(new_n862_), .C1(new_n848_), .C2(KEYINPUT59), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n861_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT124), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n869_), .B(new_n861_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1341gat));
  OAI21_X1  g670(.A(G127gat), .B1(new_n855_), .B2(new_n721_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n721_), .A2(G127gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n848_), .B2(new_n873_), .ZN(G1342gat));
  INV_X1    g673(.A(new_n661_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G134gat), .B1(new_n855_), .B2(new_n875_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n365_), .A2(G134gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n848_), .B2(new_n877_), .ZN(G1343gat));
  OR2_X1    g677(.A1(new_n843_), .A2(new_n847_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n442_), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n590_), .A2(new_n560_), .A3(new_n554_), .A4(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n615_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n400_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n297_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n401_), .ZN(G1345gat));
  NOR2_X1   g685(.A1(new_n882_), .A2(new_n721_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT61), .B(G155gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n882_), .B2(new_n875_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n365_), .A2(G162gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n882_), .B2(new_n891_), .ZN(G1347gat));
  NOR2_X1   g691(.A1(new_n595_), .A2(new_n623_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n560_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n853_), .A2(new_n442_), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n634_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G169gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n898_));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n615_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n897_), .A2(new_n898_), .B1(new_n900_), .B2(new_n467_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n897_), .B2(new_n898_), .ZN(G1348gat));
  AOI21_X1  g701(.A(G176gat), .B1(new_n895_), .B2(new_n720_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n879_), .A2(new_n880_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n894_), .A2(new_n454_), .A3(new_n297_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  NOR3_X1   g705(.A1(new_n899_), .A2(new_n457_), .A3(new_n721_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n904_), .A2(new_n560_), .A3(new_n893_), .A4(new_n325_), .ZN(new_n908_));
  INV_X1    g707(.A(G183gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n908_), .B2(new_n909_), .ZN(G1350gat));
  OAI21_X1  g709(.A(G190gat), .B1(new_n899_), .B2(new_n875_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n895_), .A2(new_n458_), .A3(new_n834_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1351gat));
  NAND3_X1  g712(.A1(new_n595_), .A2(new_n554_), .A3(new_n442_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n560_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n915_), .B2(new_n914_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n879_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n615_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(new_n382_), .ZN(G1352gat));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n297_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n380_), .ZN(G1353gat));
  INV_X1    g721(.A(new_n918_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT63), .B(G211gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n923_), .A2(new_n325_), .A3(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926_));
  OAI22_X1  g725(.A1(new_n918_), .A2(new_n721_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n925_), .B2(new_n927_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1354gat));
  OR3_X1    g729(.A1(new_n918_), .A2(G218gat), .A3(new_n365_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G218gat), .B1(new_n918_), .B2(new_n875_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1355gat));
endmodule


