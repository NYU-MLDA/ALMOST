//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n585_, new_n586_, new_n587_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  XOR2_X1   g004(.A(G197gat), .B(G204gat), .Z(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(KEYINPUT21), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(KEYINPUT21), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n208_), .A2(new_n209_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT22), .B(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n217_), .B2(KEYINPUT22), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n213_), .B1(new_n216_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT85), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n222_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT86), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n226_), .B2(KEYINPUT23), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n225_), .A2(new_n229_), .A3(new_n227_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n223_), .B(new_n224_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  OR3_X1    g034(.A1(new_n226_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT83), .B1(new_n226_), .B2(KEYINPUT23), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n236_), .B(new_n237_), .C1(new_n225_), .C2(new_n227_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT25), .B(G183gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT26), .B(G190gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n239_), .A2(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n238_), .B(new_n243_), .C1(new_n242_), .C2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n235_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT87), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT87), .B1(new_n235_), .B2(new_n245_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n212_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n212_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n242_), .B1(new_n244_), .B2(KEYINPUT93), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(KEYINPUT93), .B2(new_n244_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n253_), .A2(new_n231_), .A3(new_n232_), .A4(new_n243_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT94), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n213_), .B(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n219_), .B2(new_n214_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT95), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(KEYINPUT95), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n238_), .B1(G183gat), .B2(G190gat), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n258_), .B(new_n259_), .C1(KEYINPUT96), .C2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n260_), .A2(KEYINPUT96), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n251_), .B(new_n254_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n263_), .A2(KEYINPUT20), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n250_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n248_), .A2(new_n212_), .A3(new_n249_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n254_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n212_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT20), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n271_), .A2(new_n274_), .A3(new_n267_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n205_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n205_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n267_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n250_), .A2(new_n268_), .A3(new_n264_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(KEYINPUT97), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT97), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n282_), .B(new_n267_), .C1(new_n271_), .C2(new_n274_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n278_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT27), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n277_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n281_), .A2(new_n278_), .A3(new_n283_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n287_), .B2(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT100), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT100), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n290_), .B(new_n285_), .C1(new_n287_), .C2(new_n284_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299_));
  OAI22_X1  g098(.A1(new_n296_), .A2(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n297_), .B2(new_n296_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n299_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT90), .ZN(new_n303_));
  AOI211_X1 g102(.A(new_n294_), .B(new_n295_), .C1(new_n301_), .C2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n298_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n295_), .B1(KEYINPUT1), .B2(new_n293_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n293_), .A2(KEYINPUT1), .ZN(new_n307_));
  AOI211_X1 g106(.A(new_n305_), .B(new_n296_), .C1(new_n306_), .C2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G22gat), .B(G50gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT28), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n311_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G228gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT91), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n309_), .A2(new_n310_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(new_n251_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n212_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n315_), .B(KEYINPUT91), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G78gat), .B(G106gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n314_), .B1(new_n325_), .B2(KEYINPUT92), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n322_), .B(new_n323_), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  XOR2_X1   g127(.A(G127gat), .B(G134gat), .Z(new_n329_));
  XOR2_X1   g128(.A(G113gat), .B(G120gat), .Z(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n309_), .A2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n334_), .A2(KEYINPUT4), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n340_), .B1(new_n335_), .B2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n339_), .B1(new_n342_), .B2(new_n338_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT0), .B(G57gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  XNOR2_X1  g146(.A(new_n343_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n328_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n348_), .B1(new_n353_), .B2(KEYINPUT99), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n281_), .A2(new_n283_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n351_), .B(KEYINPUT98), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n354_), .B(new_n357_), .C1(KEYINPUT99), .C2(new_n353_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n287_), .A2(new_n284_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT33), .ZN(new_n360_));
  INV_X1    g159(.A(new_n347_), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n343_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n347_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n360_), .B1(new_n343_), .B2(new_n361_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n359_), .A2(new_n362_), .A3(new_n364_), .A4(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n358_), .A2(new_n366_), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n292_), .A2(new_n350_), .B1(new_n367_), .B2(new_n328_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n248_), .A2(new_n249_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT88), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT30), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n369_), .B(new_n372_), .Z(new_n373_));
  XOR2_X1   g172(.A(G71gat), .B(G99gat), .Z(new_n374_));
  OR2_X1    g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n374_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT31), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n332_), .B2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n379_), .B2(new_n332_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G15gat), .B(G43gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n377_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n375_), .A2(new_n383_), .A3(new_n376_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n328_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n292_), .ZN(new_n391_));
  OAI22_X1  g190(.A1(new_n368_), .A2(new_n388_), .B1(new_n349_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT76), .B(G15gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G22gat), .ZN(new_n395_));
  INV_X1    g194(.A(G1gat), .ZN(new_n396_));
  INV_X1    g195(.A(G8gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT14), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G1gat), .B(G8gat), .Z(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G29gat), .B(G36gat), .Z(new_n402_));
  XOR2_X1   g201(.A(G43gat), .B(G50gat), .Z(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT79), .ZN(new_n407_));
  INV_X1    g206(.A(new_n401_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n404_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n407_), .B(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G229gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n404_), .B(KEYINPUT15), .Z(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n408_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n411_), .A3(new_n406_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n393_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G113gat), .B(G141gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G169gat), .B(G197gat), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(new_n421_), .Z(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n418_), .B1(new_n422_), .B2(new_n393_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n419_), .A2(new_n423_), .B1(new_n425_), .B2(new_n417_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G127gat), .B(G155gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT16), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G183gat), .B(G211gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT17), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT78), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G57gat), .B(G64gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT11), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT68), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT68), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(new_n437_), .A3(KEYINPUT11), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n434_), .A2(KEYINPUT11), .ZN(new_n440_));
  XOR2_X1   g239(.A(G71gat), .B(G78gat), .Z(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n436_), .A2(new_n440_), .A3(new_n441_), .A4(new_n438_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n401_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G231gat), .A2(G233gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n433_), .B1(new_n448_), .B2(KEYINPUT77), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(KEYINPUT77), .B2(new_n448_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n430_), .A2(new_n431_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(G85gat), .ZN(new_n454_));
  INV_X1    g253(.A(G92gat), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n454_), .A2(new_n455_), .A3(KEYINPUT9), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G85gat), .B(G92gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n456_), .B1(new_n458_), .B2(KEYINPUT9), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT10), .B(G99gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G99gat), .A2(G106gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT6), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(G99gat), .A3(G106gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n467_), .A3(KEYINPUT65), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n466_), .B1(G99gat), .B2(G106gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n464_), .A2(KEYINPUT6), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n459_), .A2(new_n463_), .A3(new_n468_), .A4(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n465_), .A2(new_n467_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n457_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT8), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT67), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n472_), .A2(new_n468_), .A3(new_n477_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n457_), .A2(KEYINPUT8), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(KEYINPUT66), .A3(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n470_), .A2(new_n471_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n486_));
  INV_X1    g285(.A(G99gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n462_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n474_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n458_), .B1(new_n485_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT67), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT8), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n481_), .A2(new_n484_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT66), .B1(new_n482_), .B2(new_n483_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n473_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT34), .ZN(new_n497_));
  OAI22_X1  g296(.A1(new_n495_), .A2(new_n404_), .B1(KEYINPUT35), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n498_), .B1(new_n414_), .B2(new_n495_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(KEYINPUT35), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G190gat), .B(G218gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT71), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G134gat), .B(G162gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n501_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n505_), .B(KEYINPUT36), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n501_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n510_), .B2(KEYINPUT72), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n501_), .A2(KEYINPUT72), .A3(new_n509_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT37), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(KEYINPUT73), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n501_), .A2(new_n509_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT73), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n514_), .A2(new_n508_), .A3(new_n517_), .A4(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n513_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT75), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT75), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n513_), .A2(new_n522_), .A3(new_n519_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n453_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n525_));
  INV_X1    g324(.A(new_n445_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n495_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT66), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n465_), .A2(new_n467_), .A3(KEYINPUT65), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT65), .B1(new_n465_), .B2(new_n467_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n489_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n483_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n528_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n533_), .A2(new_n484_), .A3(new_n481_), .A4(new_n492_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(new_n473_), .A3(new_n445_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n525_), .B1(new_n527_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G230gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT64), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n495_), .A2(new_n526_), .B1(new_n540_), .B2(KEYINPUT12), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n536_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n538_), .B1(new_n527_), .B2(new_n535_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G120gat), .B(G148gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT5), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G176gat), .B(G204gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n548_), .B(KEYINPUT70), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n544_), .A2(new_n552_), .ZN(new_n553_));
  OR3_X1    g352(.A1(new_n550_), .A2(new_n553_), .A3(KEYINPUT13), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT13), .B1(new_n550_), .B2(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n392_), .A2(new_n426_), .A3(new_n524_), .A4(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n348_), .B(KEYINPUT101), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n557_), .A2(G1gat), .A3(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n514_), .A2(new_n508_), .A3(new_n517_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n392_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n556_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n426_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n453_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(G1gat), .B1(new_n568_), .B2(new_n348_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n560_), .A2(new_n561_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT103), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n570_), .A2(new_n571_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n562_), .B(new_n569_), .C1(new_n573_), .C2(new_n574_), .ZN(G1324gat));
  NOR3_X1   g374(.A1(new_n557_), .A2(G8gat), .A3(new_n292_), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT104), .Z(new_n577_));
  OAI21_X1  g376(.A(G8gat), .B1(new_n568_), .B2(new_n292_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT39), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT40), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(G1325gat));
  OAI21_X1  g383(.A(G15gat), .B1(new_n568_), .B2(new_n387_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT41), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n557_), .A2(G15gat), .A3(new_n387_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(new_n587_), .ZN(G1326gat));
  OAI21_X1  g387(.A(G22gat), .B1(new_n568_), .B2(new_n328_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n328_), .A2(G22gat), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n591_), .B1(new_n557_), .B2(new_n592_), .ZN(G1327gat));
  NAND2_X1  g392(.A1(new_n521_), .A2(new_n523_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n292_), .A2(new_n350_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n367_), .A2(new_n328_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n388_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n390_), .A2(new_n292_), .A3(new_n348_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n595_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT43), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT43), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n392_), .A2(new_n602_), .A3(new_n595_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n565_), .A2(new_n566_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n453_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT44), .B1(new_n604_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT44), .ZN(new_n609_));
  AOI211_X1 g408(.A(new_n609_), .B(new_n606_), .C1(new_n601_), .C2(new_n603_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n608_), .A2(new_n610_), .A3(new_n559_), .ZN(new_n611_));
  INV_X1    g410(.A(G29gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n453_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n563_), .A2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n614_), .A2(new_n556_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n392_), .A2(new_n426_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n349_), .A2(new_n612_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT106), .ZN(new_n618_));
  OAI22_X1  g417(.A1(new_n611_), .A2(new_n612_), .B1(new_n616_), .B2(new_n618_), .ZN(G1328gat));
  NAND2_X1  g418(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT108), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT46), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(G36gat), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n608_), .A2(new_n610_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n292_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n292_), .A2(G36gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OR3_X1    g428(.A1(new_n616_), .A2(KEYINPUT107), .A3(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT107), .B1(new_n616_), .B2(new_n629_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT45), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n630_), .A2(KEYINPUT45), .A3(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n620_), .B(new_n623_), .C1(new_n627_), .C2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n608_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n604_), .A2(KEYINPUT44), .A3(new_n607_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n626_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G36gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n635_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT45), .B1(new_n630_), .B2(new_n631_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n641_), .A2(new_n644_), .A3(new_n621_), .A4(new_n622_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n637_), .A2(new_n645_), .ZN(G1329gat));
  INV_X1    g445(.A(new_n616_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G43gat), .B1(new_n647_), .B2(new_n388_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n388_), .A2(G43gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n625_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g450(.A(G50gat), .B1(new_n647_), .B2(new_n389_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n389_), .A2(G50gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n625_), .B2(new_n653_), .ZN(G1331gat));
  NOR2_X1   g453(.A1(new_n556_), .A2(new_n426_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n564_), .A2(new_n613_), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G57gat), .B1(new_n656_), .B2(new_n348_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n392_), .A2(new_n655_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n524_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n559_), .A2(G57gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(G1332gat));
  OAI21_X1  g460(.A(G64gat), .B1(new_n656_), .B2(new_n292_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT48), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n292_), .A2(G64gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n659_), .B2(new_n664_), .ZN(G1333gat));
  OAI21_X1  g464(.A(G71gat), .B1(new_n656_), .B2(new_n387_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT49), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n387_), .A2(G71gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n659_), .B2(new_n668_), .ZN(G1334gat));
  OAI21_X1  g468(.A(G78gat), .B1(new_n656_), .B2(new_n328_), .ZN(new_n670_));
  XOR2_X1   g469(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n328_), .A2(G78gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n659_), .B2(new_n673_), .ZN(G1335gat));
  NAND3_X1  g473(.A1(new_n601_), .A2(KEYINPUT110), .A3(new_n603_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT110), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n604_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n675_), .A2(new_n453_), .A3(new_n655_), .A4(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G85gat), .B1(new_n678_), .B2(new_n348_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n658_), .A2(new_n614_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n454_), .A3(new_n558_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(G1336gat));
  OAI21_X1  g482(.A(G92gat), .B1(new_n678_), .B2(new_n292_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(new_n455_), .A3(new_n626_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT111), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n688_), .A3(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1337gat));
  OAI21_X1  g489(.A(G99gat), .B1(new_n678_), .B2(new_n387_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n681_), .A2(new_n388_), .A3(new_n461_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT51), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT51), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n691_), .A2(new_n695_), .A3(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1338gat));
  NAND3_X1  g496(.A1(new_n681_), .A2(new_n462_), .A3(new_n389_), .ZN(new_n698_));
  NOR4_X1   g497(.A1(new_n556_), .A2(new_n426_), .A3(new_n328_), .A4(new_n613_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n462_), .B1(new_n604_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT52), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n700_), .A2(new_n701_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n698_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT53), .ZN(G1339gat));
  XOR2_X1   g504(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n706_));
  AND3_X1   g505(.A1(new_n513_), .A2(new_n522_), .A3(new_n519_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n522_), .B1(new_n513_), .B2(new_n519_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n613_), .B(new_n556_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n706_), .B1(new_n709_), .B2(new_n426_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT54), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n711_), .A2(KEYINPUT112), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n524_), .A2(new_n566_), .A3(new_n556_), .A4(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n710_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n413_), .A2(new_n422_), .A3(new_n416_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n411_), .B1(new_n415_), .B2(new_n406_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n410_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(new_n411_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n716_), .B1(new_n719_), .B2(new_n422_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(new_n550_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT118), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n539_), .B1(new_n536_), .B2(new_n541_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n525_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n534_), .A2(new_n473_), .A3(new_n445_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n445_), .B1(new_n534_), .B2(new_n473_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n540_), .A2(KEYINPUT12), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n527_), .A2(new_n728_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n727_), .A2(KEYINPUT55), .A3(new_n538_), .A4(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n723_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n727_), .A2(new_n538_), .A3(new_n729_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n731_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT113), .B1(new_n542_), .B2(KEYINPUT55), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(KEYINPUT114), .A3(new_n731_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n552_), .B1(new_n739_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n722_), .B1(new_n744_), .B2(KEYINPUT56), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT114), .B1(new_n742_), .B2(new_n731_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n723_), .A2(new_n730_), .ZN(new_n747_));
  AOI211_X1 g546(.A(new_n738_), .B(new_n747_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n551_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(KEYINPUT118), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n745_), .A2(new_n751_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT56), .B(new_n551_), .C1(new_n746_), .C2(new_n748_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n744_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n721_), .B1(new_n752_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI211_X1 g559(.A(KEYINPUT58), .B(new_n721_), .C1(new_n752_), .C2(new_n757_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n595_), .A3(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT57), .ZN(new_n763_));
  INV_X1    g562(.A(new_n563_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n750_), .B1(new_n744_), .B2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n749_), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n426_), .A2(new_n549_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n550_), .A2(new_n553_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n720_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n763_), .B(new_n764_), .C1(new_n770_), .C2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n764_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(KEYINPUT57), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n739_), .A2(new_n743_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n765_), .B1(new_n779_), .B2(new_n551_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n768_), .B1(new_n780_), .B2(KEYINPUT56), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n772_), .B1(new_n781_), .B2(new_n766_), .ZN(new_n782_));
  OAI211_X1 g581(.A(KEYINPUT116), .B(new_n763_), .C1(new_n782_), .C2(new_n764_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n762_), .A2(new_n775_), .A3(new_n778_), .A4(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n715_), .B1(new_n784_), .B2(new_n453_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n391_), .A2(new_n559_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(G113gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n426_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT59), .B1(new_n785_), .B2(new_n787_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n793_));
  AOI21_X1  g592(.A(new_n594_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n774_), .B1(new_n794_), .B2(new_n761_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n763_), .B1(new_n782_), .B2(new_n764_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n613_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n786_), .B(new_n793_), .C1(new_n797_), .C2(new_n715_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n791_), .A2(new_n792_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n792_), .B1(new_n791_), .B2(new_n798_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n799_), .A2(new_n800_), .A3(new_n566_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n790_), .B1(new_n801_), .B2(new_n789_), .ZN(G1340gat));
  INV_X1    g601(.A(KEYINPUT60), .ZN(new_n803_));
  AOI21_X1  g602(.A(G120gat), .B1(new_n565_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n803_), .B2(G120gat), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n788_), .A2(new_n805_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(KEYINPUT121), .Z(new_n807_));
  NAND3_X1  g606(.A1(new_n791_), .A2(new_n565_), .A3(new_n798_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(G120gat), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(G1341gat));
  INV_X1    g609(.A(G127gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n788_), .A2(new_n811_), .A3(new_n613_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n799_), .A2(new_n800_), .A3(new_n453_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n811_), .ZN(G1342gat));
  INV_X1    g613(.A(G134gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n788_), .A2(new_n815_), .A3(new_n764_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n799_), .A2(new_n800_), .A3(new_n594_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n815_), .ZN(G1343gat));
  INV_X1    g617(.A(new_n785_), .ZN(new_n819_));
  NOR4_X1   g618(.A1(new_n626_), .A2(new_n328_), .A3(new_n388_), .A4(new_n559_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(new_n566_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT122), .B(G141gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1344gat));
  NOR2_X1   g623(.A1(new_n821_), .A2(new_n556_), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n825_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g625(.A1(new_n821_), .A2(new_n453_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT61), .B(G155gat), .Z(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(G1346gat));
  NAND2_X1  g628(.A1(new_n595_), .A2(G162gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT124), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n819_), .A2(new_n820_), .A3(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n778_), .A2(new_n783_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n613_), .B1(new_n833_), .B2(new_n795_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n764_), .B(new_n820_), .C1(new_n834_), .C2(new_n715_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n836_));
  INV_X1    g635(.A(G162gat), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n832_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT125), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n842_), .B(new_n832_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1347gat));
  OR2_X1    g643(.A1(new_n797_), .A2(new_n715_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n292_), .A2(new_n387_), .A3(new_n558_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n328_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(G169gat), .B1(new_n847_), .B2(new_n566_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n845_), .A2(new_n328_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n851_), .A2(new_n426_), .A3(new_n214_), .A4(new_n846_), .ZN(new_n852_));
  OAI211_X1 g651(.A(KEYINPUT62), .B(G169gat), .C1(new_n847_), .C2(new_n566_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(new_n852_), .A3(new_n853_), .ZN(G1348gat));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n565_), .A3(new_n846_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n785_), .A2(new_n389_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n846_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n857_), .A2(new_n219_), .A3(new_n556_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n855_), .A2(new_n219_), .B1(new_n856_), .B2(new_n858_), .ZN(G1349gat));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n453_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G183gat), .B1(new_n856_), .B2(new_n860_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n857_), .A2(new_n239_), .A3(new_n453_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n851_), .B2(new_n862_), .ZN(G1350gat));
  OAI21_X1  g662(.A(G190gat), .B1(new_n847_), .B2(new_n594_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n764_), .A2(new_n240_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n847_), .B2(new_n865_), .ZN(G1351gat));
  NAND2_X1  g665(.A1(new_n387_), .A2(new_n350_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT126), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n785_), .A2(new_n292_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n426_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n565_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g672(.A(KEYINPUT63), .B(G211gat), .C1(new_n869_), .C2(new_n613_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n869_), .A2(new_n613_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT63), .B(G211gat), .Z(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(G1354gat));
  AOI21_X1  g676(.A(G218gat), .B1(new_n869_), .B2(new_n764_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n595_), .A2(G218gat), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT127), .Z(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n869_), .B2(new_n880_), .ZN(G1355gat));
endmodule


