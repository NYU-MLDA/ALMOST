//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_;
  OR3_X1    g000(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT23), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n207_), .B2(KEYINPUT23), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G183gat), .ZN(new_n212_));
  INV_X1    g011(.A(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n204_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT91), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G218gat), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n218_), .A2(G211gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(G211gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT86), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G211gat), .B(G218gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT86), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G197gat), .ZN(new_n225_));
  INV_X1    g024(.A(G204gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n227_), .A2(KEYINPUT21), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n221_), .A2(new_n224_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT87), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n224_), .A2(new_n221_), .A3(new_n229_), .A4(KEYINPUT87), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n227_), .A2(new_n228_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(KEYINPUT21), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n227_), .A2(KEYINPUT21), .A3(new_n228_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n236_), .A2(new_n222_), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n232_), .A2(new_n233_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n212_), .A2(KEYINPUT25), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G183gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n213_), .A2(KEYINPUT26), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT26), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G190gat), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n239_), .A2(new_n241_), .A3(new_n242_), .A4(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT24), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n207_), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT76), .B1(new_n207_), .B2(KEYINPUT23), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n206_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n246_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(KEYINPUT24), .A3(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n249_), .A2(new_n252_), .A3(KEYINPUT90), .A4(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT90), .ZN(new_n257_));
  INV_X1    g056(.A(new_n206_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n251_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n207_), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n245_), .A2(new_n255_), .A3(new_n248_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n257_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n256_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n217_), .A2(new_n238_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT20), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n232_), .A2(new_n233_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n235_), .A2(new_n237_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n204_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n214_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n270_), .B1(new_n261_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n211_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n272_), .B1(new_n262_), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n266_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT19), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n265_), .A2(new_n275_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT92), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n211_), .A2(new_n214_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n216_), .B1(new_n281_), .B2(new_n270_), .ZN(new_n282_));
  AOI211_X1 g081(.A(KEYINPUT91), .B(new_n204_), .C1(new_n211_), .C2(new_n214_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n256_), .A2(new_n263_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n269_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n204_), .B1(new_n252_), .B2(new_n214_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n262_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(new_n211_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n266_), .B1(new_n238_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n280_), .B1(new_n291_), .B2(new_n277_), .ZN(new_n292_));
  AOI211_X1 g091(.A(KEYINPUT92), .B(new_n278_), .C1(new_n286_), .C2(new_n290_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n279_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT18), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT32), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT98), .ZN(new_n301_));
  INV_X1    g100(.A(new_n275_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n261_), .A2(new_n262_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n269_), .A2(new_n303_), .A3(new_n215_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n277_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(new_n277_), .B2(new_n291_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n300_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n295_), .A2(new_n301_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT95), .ZN(new_n309_));
  XOR2_X1   g108(.A(G141gat), .B(G148gat), .Z(new_n310_));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(G155gat), .A3(G162gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n312_), .B(KEYINPUT82), .Z(new_n313_));
  INV_X1    g112(.A(KEYINPUT81), .ZN(new_n314_));
  INV_X1    g113(.A(G155gat), .ZN(new_n315_));
  INV_X1    g114(.A(G162gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n319_), .B1(new_n311_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n310_), .B1(new_n313_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT84), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n320_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT83), .ZN(new_n326_));
  OR3_X1    g125(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n323_), .B(new_n324_), .C1(new_n326_), .C2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n328_), .A2(new_n329_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT83), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n325_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n325_), .A2(new_n334_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n333_), .B(new_n327_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n323_), .B1(new_n337_), .B2(new_n324_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n322_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G127gat), .B(G134gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n342_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n344_), .B(new_n322_), .C1(new_n332_), .C2(new_n338_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(KEYINPUT4), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT94), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n343_), .A2(new_n345_), .A3(KEYINPUT94), .A4(KEYINPUT4), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n343_), .B2(KEYINPUT4), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n309_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n343_), .A2(new_n345_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(new_n352_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n353_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(KEYINPUT95), .ZN(new_n358_));
  XOR2_X1   g157(.A(KEYINPUT96), .B(KEYINPUT0), .Z(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT97), .ZN(new_n360_));
  XOR2_X1   g159(.A(G1gat), .B(G29gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n354_), .A2(new_n358_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n308_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT33), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n354_), .A2(new_n358_), .A3(KEYINPUT33), .A4(new_n365_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n238_), .B1(new_n217_), .B2(new_n264_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT20), .B1(new_n269_), .B2(new_n274_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n277_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT92), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n291_), .A2(new_n280_), .A3(new_n277_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n299_), .B1(new_n379_), .B2(new_n279_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n299_), .B(new_n279_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT93), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n299_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n294_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n381_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n351_), .B1(new_n343_), .B2(KEYINPUT4), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n364_), .B1(new_n355_), .B2(new_n351_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n383_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n369_), .B1(new_n373_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n238_), .B1(new_n339_), .B2(KEYINPUT29), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT88), .B1(G228gat), .B2(G233gat), .ZN(new_n396_));
  AND3_X1   g195(.A1(KEYINPUT88), .A2(G228gat), .A3(G233gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT89), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n400_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n398_), .B(new_n404_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G22gat), .B(G50gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT28), .ZN(new_n408_));
  INV_X1    g207(.A(new_n339_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n339_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n407_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n411_), .A2(new_n412_), .A3(new_n407_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n399_), .A2(new_n402_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n403_), .A2(new_n405_), .A3(new_n416_), .A4(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT85), .B1(new_n414_), .B2(new_n415_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n415_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n413_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n405_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n419_), .B(new_n422_), .C1(new_n401_), .C2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n394_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT99), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n418_), .A2(new_n424_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n385_), .A2(new_n381_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n391_), .B1(new_n429_), .B2(KEYINPUT93), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n430_), .A2(new_n387_), .A3(new_n371_), .A4(new_n372_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n428_), .B1(new_n431_), .B2(new_n369_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT99), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n382_), .A2(KEYINPUT100), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT100), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n381_), .A2(new_n437_), .B1(new_n306_), .B2(new_n384_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n435_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n429_), .A2(KEYINPUT27), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n367_), .A2(new_n368_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n428_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n427_), .A2(new_n434_), .A3(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G71gat), .B(G99gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT77), .B(G43gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  XNOR2_X1  g246(.A(new_n289_), .B(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G227gat), .A2(G233gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n449_), .B(G15gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT30), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n451_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT79), .B1(new_n454_), .B2(KEYINPUT78), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n342_), .B(KEYINPUT31), .Z(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n454_), .B2(KEYINPUT78), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT78), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT79), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n452_), .A2(new_n458_), .A3(new_n459_), .A4(new_n453_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n455_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n457_), .B1(new_n455_), .B2(new_n460_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n463_), .B(KEYINPUT80), .Z(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT101), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n425_), .B1(new_n440_), .B2(new_n439_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n442_), .A2(new_n463_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n442_), .A2(new_n463_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n470_), .A2(new_n441_), .A3(KEYINPUT101), .A4(new_n425_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n444_), .A2(new_n465_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G29gat), .B(G36gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT68), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G43gat), .B(G50gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n473_), .A2(KEYINPUT68), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(KEYINPUT68), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n475_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT15), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484_));
  INV_X1    g283(.A(G1gat), .ZN(new_n485_));
  INV_X1    g284(.A(G8gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G1gat), .B(G8gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n477_), .A2(KEYINPUT15), .A3(new_n480_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n483_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT73), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n483_), .A2(KEYINPUT73), .A3(new_n490_), .A4(new_n491_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n490_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n477_), .A2(KEYINPUT72), .A3(new_n480_), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT72), .B1(new_n477_), .B2(new_n480_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G229gat), .A2(G233gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n498_), .A2(new_n499_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n490_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n501_), .B1(new_n504_), .B2(new_n500_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n502_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n500_), .A2(new_n501_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n513_), .B2(new_n505_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n514_), .A3(KEYINPUT74), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT74), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n516_), .B(new_n511_), .C1(new_n513_), .C2(new_n505_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n472_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT6), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT65), .ZN(new_n522_));
  INV_X1    g321(.A(G99gat), .ZN(new_n523_));
  INV_X1    g322(.A(G106gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT7), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n522_), .A2(new_n527_), .A3(new_n523_), .A4(new_n524_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n521_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G85gat), .B(G92gat), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT8), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n536_));
  XOR2_X1   g335(.A(G71gat), .B(G78gat), .Z(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n536_), .A2(new_n537_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n529_), .A2(KEYINPUT8), .A3(new_n530_), .ZN(new_n541_));
  INV_X1    g340(.A(G85gat), .ZN(new_n542_));
  INV_X1    g341(.A(G92gat), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n542_), .A2(new_n543_), .A3(KEYINPUT9), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n530_), .B2(KEYINPUT9), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT64), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT10), .B(G99gat), .Z(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n547_), .B2(new_n524_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT10), .B(G99gat), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n549_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n521_), .B(new_n545_), .C1(new_n548_), .C2(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n533_), .A2(new_n540_), .A3(new_n541_), .A4(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n533_), .A2(new_n541_), .A3(new_n551_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n556_));
  INV_X1    g355(.A(new_n540_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n556_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n554_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(new_n557_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n561_), .A2(new_n552_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n553_), .B2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G120gat), .B(G148gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G176gat), .B(G204gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n563_), .B(new_n568_), .Z(new_n569_));
  INV_X1    g368(.A(KEYINPUT13), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n570_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT67), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n490_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n557_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n578_), .A2(KEYINPUT71), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT16), .ZN(new_n581_));
  XOR2_X1   g380(.A(G183gat), .B(G211gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n578_), .A2(new_n583_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n584_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n483_), .A2(new_n555_), .A3(new_n491_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n481_), .A2(new_n541_), .A3(new_n551_), .A4(new_n533_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT35), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n596_), .A2(KEYINPUT35), .A3(new_n594_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(KEYINPUT35), .B2(new_n594_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT36), .ZN(new_n602_));
  OR3_X1    g401(.A1(new_n597_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(KEYINPUT36), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n602_), .B(new_n604_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(KEYINPUT69), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n519_), .A2(new_n575_), .A3(new_n590_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  INV_X1    g410(.A(new_n442_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n485_), .ZN(new_n613_));
  OR3_X1    g412(.A1(new_n610_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n603_), .A2(new_n605_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT102), .Z(new_n616_));
  NOR2_X1   g415(.A1(new_n472_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n573_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(new_n518_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n589_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n442_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n611_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n614_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT103), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(G1324gat));
  OR3_X1    g426(.A1(new_n610_), .A2(G8gat), .A3(new_n441_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G8gat), .B1(new_n622_), .B2(new_n441_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(KEYINPUT39), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(KEYINPUT39), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n628_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT40), .B(new_n628_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n622_), .B2(new_n465_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT41), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n610_), .A2(G15gat), .A3(new_n465_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1326gat));
  XNOR2_X1  g439(.A(new_n428_), .B(KEYINPUT104), .ZN(new_n641_));
  OAI21_X1  g440(.A(G22gat), .B1(new_n622_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT42), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n641_), .A2(G22gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n643_), .B1(new_n610_), .B2(new_n644_), .ZN(G1327gat));
  INV_X1    g444(.A(new_n615_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n589_), .A2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT106), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n519_), .A2(new_n573_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n612_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n620_), .A2(new_n590_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n443_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n654_));
  AOI211_X1 g453(.A(KEYINPUT99), .B(new_n428_), .C1(new_n431_), .C2(new_n369_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n465_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n471_), .A2(new_n469_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n653_), .B1(new_n658_), .B2(new_n608_), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT43), .B(new_n609_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT44), .B(new_n652_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n652_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT43), .B1(new_n472_), .B2(new_n609_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n658_), .A2(new_n653_), .A3(new_n608_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n612_), .A2(G29gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n651_), .B1(new_n668_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(new_n441_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n661_), .B(new_n671_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G36gat), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n441_), .A2(KEYINPUT107), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n441_), .A2(KEYINPUT107), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  OR3_X1    g477(.A1(new_n649_), .A2(KEYINPUT45), .A3(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT45), .B1(new_n649_), .B2(new_n678_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n673_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n673_), .A2(new_n681_), .A3(KEYINPUT46), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1329gat));
  XNOR2_X1  g485(.A(KEYINPUT108), .B(G43gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(new_n649_), .B2(new_n465_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n463_), .A2(G43gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n667_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g490(.A(new_n641_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G50gat), .B1(new_n650_), .B2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n428_), .A2(G50gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n668_), .B2(new_n694_), .ZN(G1331gat));
  INV_X1    g494(.A(new_n518_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n472_), .A2(new_n696_), .ZN(new_n697_));
  AND4_X1   g496(.A1(new_n618_), .A2(new_n697_), .A3(new_n590_), .A4(new_n609_), .ZN(new_n698_));
  INV_X1    g497(.A(G57gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n612_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n589_), .A2(new_n696_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n617_), .A2(new_n574_), .A3(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n442_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(G1332gat));
  OAI21_X1  g503(.A(G64gat), .B1(new_n702_), .B2(new_n677_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT48), .ZN(new_n706_));
  INV_X1    g505(.A(G64gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n698_), .A2(new_n707_), .A3(new_n676_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1333gat));
  OAI21_X1  g508(.A(G71gat), .B1(new_n702_), .B2(new_n465_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT49), .ZN(new_n711_));
  INV_X1    g510(.A(G71gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n698_), .A2(new_n712_), .A3(new_n464_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1334gat));
  OAI21_X1  g513(.A(G78gat), .B1(new_n702_), .B2(new_n641_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT50), .ZN(new_n716_));
  INV_X1    g515(.A(G78gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n698_), .A2(new_n717_), .A3(new_n692_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1335gat));
  NOR3_X1   g518(.A1(new_n590_), .A2(new_n573_), .A3(new_n696_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G85gat), .B1(new_n723_), .B2(new_n442_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n697_), .A2(new_n574_), .A3(new_n648_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n542_), .A3(new_n612_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1336gat));
  OAI21_X1  g526(.A(G92gat), .B1(new_n723_), .B2(new_n677_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n543_), .A3(new_n671_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1337gat));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n463_), .A3(new_n547_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n464_), .B(new_n720_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(G99gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G99gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT51), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n738_), .B(new_n731_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1338gat));
  NAND3_X1  g539(.A1(new_n725_), .A2(new_n524_), .A3(new_n428_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n428_), .B(new_n720_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(G106gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(G106gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n741_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  INV_X1    g549(.A(G113gat), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n701_), .A2(new_n573_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n609_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(new_n609_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n560_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n561_), .A2(KEYINPUT12), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n763_), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(new_n554_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n760_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n553_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n552_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n768_));
  AOI22_X1  g567(.A1(new_n766_), .A2(new_n767_), .B1(new_n560_), .B2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n765_), .A2(KEYINPUT112), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n568_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT112), .B1(new_n765_), .B2(new_n769_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n563_), .A2(new_n568_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n504_), .A2(new_n500_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n509_), .B1(new_n775_), .B2(new_n501_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n496_), .A2(G229gat), .A3(G233gat), .A4(new_n500_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n774_), .A2(new_n510_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n765_), .A2(new_n769_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n568_), .A4(new_n770_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n773_), .A2(new_n779_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(KEYINPUT58), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n787_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n773_), .A2(new_n784_), .A3(new_n789_), .A4(new_n779_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n608_), .A3(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT116), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n778_), .A2(new_n510_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n569_), .A2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(KEYINPUT113), .A2(KEYINPUT56), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n782_), .A2(new_n568_), .A3(new_n770_), .A4(new_n795_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n515_), .A2(new_n517_), .A3(new_n774_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n797_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n794_), .B1(new_n800_), .B2(KEYINPUT114), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n797_), .A2(new_n798_), .A3(new_n799_), .A4(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n646_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n804_), .A2(KEYINPUT57), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n806_), .B(new_n646_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n792_), .A2(new_n805_), .A3(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n757_), .B1(new_n809_), .B2(new_n590_), .ZN(new_n810_));
  NOR4_X1   g609(.A1(new_n467_), .A2(new_n461_), .A3(new_n462_), .A4(new_n442_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n751_), .B1(new_n812_), .B2(new_n518_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n518_), .A2(new_n751_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n791_), .B1(new_n804_), .B2(KEYINPUT57), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n589_), .B1(new_n817_), .B2(new_n807_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT118), .B(new_n589_), .C1(new_n817_), .C2(new_n807_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n757_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n811_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n812_), .ZN(new_n826_));
  OAI221_X1 g625(.A(new_n816_), .B1(new_n823_), .B2(new_n825_), .C1(new_n826_), .C2(new_n824_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n813_), .A2(new_n814_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n815_), .A2(new_n827_), .A3(new_n828_), .ZN(G1340gat));
  INV_X1    g628(.A(G120gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n826_), .B(new_n831_), .C1(KEYINPUT60), .C2(new_n830_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n823_), .A2(new_n825_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n824_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n833_), .A2(new_n575_), .A3(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n832_), .B1(new_n835_), .B2(new_n830_), .ZN(G1341gat));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n826_), .A2(new_n837_), .A3(new_n590_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n833_), .A2(new_n589_), .A3(new_n834_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n837_), .ZN(G1342gat));
  INV_X1    g639(.A(G134gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n826_), .A2(new_n841_), .A3(new_n616_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n833_), .A2(new_n609_), .A3(new_n834_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n841_), .ZN(G1343gat));
  NAND2_X1  g643(.A1(new_n465_), .A2(new_n428_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n845_), .A2(new_n676_), .A3(new_n442_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n810_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n696_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n574_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(new_n853_), .A3(new_n590_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT119), .B1(new_n847_), .B2(new_n589_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1346gat));
  NOR2_X1   g658(.A1(new_n847_), .A2(new_n609_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n316_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n616_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n847_), .A2(G162gat), .A3(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT120), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n848_), .A2(new_n316_), .A3(new_n616_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n865_), .B(new_n866_), .C1(new_n316_), .C2(new_n860_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(G1347gat));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n465_), .A2(new_n612_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n676_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n692_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n822_), .A2(new_n869_), .A3(new_n696_), .A4(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G169gat), .ZN(new_n874_));
  INV_X1    g673(.A(new_n872_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n756_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n821_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n869_), .B1(new_n877_), .B2(new_n696_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT62), .B1(new_n874_), .B2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n822_), .A2(new_n696_), .A3(new_n872_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT121), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(G169gat), .A4(new_n873_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT22), .B(G169gat), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n696_), .A2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT122), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n877_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n888_), .ZN(G1348gat));
  AOI21_X1  g688(.A(G176gat), .B1(new_n877_), .B2(new_n618_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n810_), .A2(new_n425_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n676_), .A2(G176gat), .A3(new_n574_), .A4(new_n870_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894_));
  OR3_X1    g693(.A1(new_n890_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n890_), .B2(new_n893_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1349gat));
  INV_X1    g696(.A(new_n877_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n239_), .A2(new_n241_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(new_n589_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n891_), .A2(new_n589_), .A3(new_n871_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(G183gat), .B1(new_n901_), .B2(new_n902_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n900_), .B1(new_n903_), .B2(new_n904_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n898_), .B2(new_n609_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n877_), .A2(new_n242_), .A3(new_n244_), .A4(new_n616_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1351gat));
  OR3_X1    g707(.A1(new_n845_), .A2(KEYINPUT125), .A3(new_n612_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT125), .B1(new_n845_), .B2(new_n612_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n909_), .A2(new_n676_), .A3(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n810_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n518_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(new_n225_), .ZN(G1352gat));
  NOR2_X1   g713(.A1(new_n912_), .A2(new_n575_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(new_n226_), .ZN(G1353gat));
  OAI22_X1  g715(.A1(new_n912_), .A2(new_n589_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT63), .B(G211gat), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n810_), .A2(new_n590_), .A3(new_n911_), .A4(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(new_n918_), .A3(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n918_), .B1(new_n917_), .B2(new_n920_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1354gat));
  NOR3_X1   g723(.A1(new_n912_), .A2(new_n218_), .A3(new_n609_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n912_), .A2(KEYINPUT127), .A3(new_n862_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(G218gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT127), .B1(new_n912_), .B2(new_n862_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n925_), .B1(new_n927_), .B2(new_n928_), .ZN(G1355gat));
endmodule


