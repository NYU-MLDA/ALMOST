//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G106gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G85gat), .ZN(new_n220_));
  INV_X1    g019(.A(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(KEYINPUT9), .A3(new_n213_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n212_), .A2(new_n214_), .A3(new_n219_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n213_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NOR3_X1   g026(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AOI211_X1 g028(.A(KEYINPUT8), .B(new_n225_), .C1(new_n229_), .C2(new_n219_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT7), .ZN(new_n232_));
  INV_X1    g031(.A(G99gat), .ZN(new_n233_));
  INV_X1    g032(.A(G106gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n217_), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n226_), .B(new_n235_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n225_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n231_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n224_), .B1(new_n230_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(KEYINPUT65), .B(new_n224_), .C1(new_n230_), .C2(new_n240_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n208_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n245_), .A2(KEYINPUT12), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(new_n208_), .A3(new_n244_), .ZN(new_n247_));
  INV_X1    g046(.A(G230gat), .ZN(new_n248_));
  INV_X1    g047(.A(G233gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n208_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n241_), .A2(new_n254_), .A3(KEYINPUT12), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n246_), .A2(new_n253_), .A3(KEYINPUT67), .A4(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n245_), .B2(KEYINPUT12), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(new_n252_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n243_), .A2(new_n244_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n254_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n251_), .B1(new_n262_), .B2(new_n247_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT66), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G120gat), .B(G148gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G176gat), .B(G204gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n260_), .A2(new_n264_), .A3(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n271_), .A2(KEYINPUT13), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT13), .B1(new_n271_), .B2(new_n273_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(KEYINPUT69), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(KEYINPUT69), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G8gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT76), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G15gat), .ZN(new_n283_));
  INV_X1    g082(.A(G22gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G15gat), .A2(G22gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G1gat), .A2(G8gat), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n285_), .A2(new_n286_), .B1(KEYINPUT14), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n282_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G29gat), .B(G36gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G43gat), .B(G50gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n289_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G229gat), .A2(G233gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n289_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n292_), .B(KEYINPUT15), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n289_), .A2(new_n292_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n294_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G113gat), .B(G141gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G169gat), .B(G197gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  NOR2_X1   g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT81), .ZN(new_n309_));
  INV_X1    g108(.A(new_n307_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n310_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n308_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n309_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT82), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(KEYINPUT82), .A3(new_n314_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n279_), .A2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G1gat), .B(G29gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT101), .B(G85gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT0), .B(G57gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G225gat), .A2(G233gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(G155gat), .B(G162gat), .Z(new_n327_));
  OR2_X1    g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT92), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n328_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT2), .Z(new_n333_));
  OAI21_X1  g132(.A(new_n327_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT1), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(G155gat), .A3(G162gat), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(new_n338_), .C1(G155gat), .C2(G162gat), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n328_), .A2(new_n332_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n339_), .A2(KEYINPUT91), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT91), .B1(new_n339_), .B2(new_n340_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n334_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G127gat), .B(G134gat), .Z(new_n344_));
  XOR2_X1   g143(.A(G113gat), .B(G120gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n346_), .B(new_n334_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT4), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n343_), .A2(new_n351_), .A3(new_n347_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n326_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n326_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n325_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT33), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT33), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n358_), .B(new_n325_), .C1(new_n353_), .C2(new_n355_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n350_), .A2(new_n326_), .A3(new_n352_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT102), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n348_), .A2(new_n349_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n325_), .B1(new_n362_), .B2(new_n354_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT102), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n350_), .A2(new_n364_), .A3(new_n326_), .A4(new_n352_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n357_), .A2(new_n359_), .B1(new_n361_), .B2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G8gat), .B(G36gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT18), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT19), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G183gat), .ZN(new_n376_));
  INV_X1    g175(.A(G190gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT23), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(G183gat), .A3(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n381_), .B1(G183gat), .B2(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT22), .B(G169gat), .ZN(new_n385_));
  INV_X1    g184(.A(G176gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n378_), .A2(KEYINPUT88), .A3(new_n380_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n390_), .B(KEYINPUT23), .C1(new_n376_), .C2(new_n377_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  OR3_X1    g191(.A1(KEYINPUT85), .A2(G169gat), .A3(G176gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(KEYINPUT24), .A3(new_n383_), .A4(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396_));
  INV_X1    g195(.A(new_n394_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(KEYINPUT85), .A2(G169gat), .A3(G176gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G190gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT25), .B(G183gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n395_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n388_), .B1(new_n392_), .B2(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(G197gat), .A2(G204gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G197gat), .A2(G204gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT21), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(KEYINPUT21), .A3(new_n406_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G211gat), .B(G218gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n410_), .A2(new_n411_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n404_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT99), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT99), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n404_), .A2(new_n417_), .A3(new_n414_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT83), .B(G183gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(new_n376_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT25), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  OR3_X1    g222(.A1(new_n376_), .A2(KEYINPUT84), .A3(KEYINPUT25), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n400_), .A3(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n425_), .A2(new_n399_), .A3(new_n395_), .A4(new_n381_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n414_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n420_), .A2(new_n377_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G169gat), .ZN(new_n431_));
  INV_X1    g230(.A(G169gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(KEYINPUT86), .A3(KEYINPUT22), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n433_), .A3(new_n386_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n435_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n429_), .B(new_n383_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n426_), .A2(new_n427_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT20), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n375_), .B1(new_n419_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n374_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n404_), .B2(new_n414_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n426_), .A2(new_n438_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(new_n414_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n372_), .B1(new_n442_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n440_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n449_), .B(new_n371_), .C1(new_n450_), .C2(new_n375_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT100), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n448_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n452_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n367_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT103), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n367_), .B(KEYINPUT103), .C1(new_n453_), .C2(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n371_), .A2(KEYINPUT32), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT97), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n414_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n404_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n443_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT105), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n463_), .A2(new_n464_), .B1(new_n446_), .B2(new_n414_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n427_), .A2(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n414_), .A2(KEYINPUT97), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT20), .B1(new_n468_), .B2(new_n404_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT105), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n374_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n450_), .A2(new_n375_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n459_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OR3_X1    g273(.A1(new_n353_), .A2(new_n325_), .A3(new_n355_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n356_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n459_), .B(KEYINPUT104), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n477_), .B(new_n449_), .C1(new_n375_), .C2(new_n450_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n457_), .A2(new_n458_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G78gat), .B(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n343_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT96), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n486_), .A2(new_n487_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n343_), .A2(KEYINPUT96), .A3(new_n485_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n484_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n414_), .A2(new_n484_), .ZN(new_n491_));
  AOI211_X1 g290(.A(KEYINPUT94), .B(new_n491_), .C1(new_n343_), .C2(KEYINPUT29), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n343_), .A2(KEYINPUT29), .ZN(new_n494_));
  INV_X1    g293(.A(new_n491_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n483_), .B1(new_n490_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n486_), .A2(new_n487_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n489_), .A3(new_n468_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n484_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n496_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n494_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n505_), .A3(new_n482_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n498_), .A2(new_n506_), .A3(KEYINPUT93), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT98), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT98), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n498_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n343_), .A2(KEYINPUT29), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT28), .ZN(new_n512_));
  XOR2_X1   g311(.A(G22gat), .B(G50gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n508_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n507_), .A2(new_n514_), .A3(KEYINPUT98), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n375_), .B1(new_n465_), .B2(new_n470_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n473_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n372_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n451_), .A2(KEYINPUT27), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n448_), .A2(new_n451_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT27), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n521_), .A2(new_n522_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n516_), .A2(new_n517_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n476_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n481_), .A2(new_n518_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G227gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(G71gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(new_n233_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n446_), .B(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G15gat), .B(G43gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT89), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT30), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n347_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT106), .B1(new_n528_), .B2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n516_), .A2(new_n517_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n525_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n541_), .A3(new_n527_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT106), .ZN(new_n547_));
  INV_X1    g346(.A(new_n541_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n474_), .A2(new_n479_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n543_), .B1(new_n550_), .B2(new_n458_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n518_), .A2(new_n544_), .A3(new_n476_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n547_), .B(new_n548_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n542_), .A2(new_n546_), .A3(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n320_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n208_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(new_n297_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G127gat), .B(G155gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT78), .ZN(new_n560_));
  XOR2_X1   g359(.A(G183gat), .B(G211gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n564_), .A2(new_n565_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n558_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n558_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT37), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT34), .Z(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n298_), .A2(new_n241_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n243_), .A2(new_n292_), .A3(new_n244_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n575_), .A2(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT71), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n580_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(KEYINPUT71), .A3(new_n582_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n578_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n581_), .A2(new_n578_), .A3(new_n582_), .A4(new_n579_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT36), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n573_), .B1(new_n587_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n586_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT71), .B1(new_n581_), .B2(new_n582_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n580_), .ZN(new_n598_));
  OAI211_X1 g397(.A(KEYINPUT72), .B(new_n595_), .C1(new_n598_), .C2(new_n578_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n594_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n591_), .B(KEYINPUT36), .Z(new_n601_));
  INV_X1    g400(.A(new_n588_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n601_), .B1(new_n587_), .B2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n572_), .B1(new_n600_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n583_), .A2(new_n584_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n586_), .A3(new_n579_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n577_), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT72), .B1(new_n608_), .B2(new_n595_), .ZN(new_n609_));
  AOI211_X1 g408(.A(new_n573_), .B(new_n593_), .C1(new_n607_), .C2(new_n577_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n572_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n601_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT73), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n587_), .B2(new_n602_), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT73), .B(new_n588_), .C1(new_n598_), .C2(new_n578_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n611_), .A2(new_n616_), .A3(KEYINPUT74), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT74), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT73), .B1(new_n608_), .B2(new_n588_), .ZN(new_n619_));
  AOI211_X1 g418(.A(new_n613_), .B(new_n602_), .C1(new_n607_), .C2(new_n577_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n601_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT37), .B1(new_n594_), .B2(new_n599_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n618_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n605_), .B1(new_n617_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT75), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT74), .B1(new_n611_), .B2(new_n616_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n621_), .A2(new_n618_), .A3(new_n622_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(KEYINPUT75), .A3(new_n605_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n571_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n555_), .A2(new_n631_), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n632_), .A2(G1gat), .A3(new_n527_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n621_), .A2(new_n600_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n554_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n279_), .A2(new_n315_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n571_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n527_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n633_), .A2(new_n634_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n641_), .A3(new_n642_), .ZN(G1324gat));
  XNOR2_X1  g442(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n644_));
  OAI21_X1  g443(.A(G8gat), .B1(new_n640_), .B2(new_n525_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT39), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n525_), .A2(G8gat), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n320_), .A2(new_n631_), .A3(new_n554_), .A4(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT107), .Z(new_n649_));
  AOI21_X1  g448(.A(new_n644_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n645_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n645_), .A2(new_n651_), .ZN(new_n653_));
  AND4_X1   g452(.A1(new_n649_), .A2(new_n652_), .A3(new_n653_), .A4(new_n644_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n650_), .A2(new_n654_), .ZN(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n640_), .B2(new_n548_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT41), .Z(new_n657_));
  INV_X1    g456(.A(new_n632_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n283_), .A3(new_n541_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(G1326gat));
  OAI21_X1  g459(.A(G22gat), .B1(new_n640_), .B2(new_n518_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT42), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(new_n284_), .A3(new_n543_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n636_), .A2(new_n570_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n555_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G29gat), .B1(new_n667_), .B2(new_n476_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT75), .B1(new_n629_), .B2(new_n605_), .ZN(new_n669_));
  AOI211_X1 g468(.A(new_n625_), .B(new_n604_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT109), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n626_), .A2(new_n672_), .A3(new_n630_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n554_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT43), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n669_), .A2(new_n670_), .A3(KEYINPUT43), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n554_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n638_), .A2(new_n570_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(KEYINPUT44), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n674_), .A2(KEYINPUT43), .B1(new_n554_), .B2(new_n676_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n679_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n680_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n476_), .A2(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n668_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  NAND3_X1  g486(.A1(new_n680_), .A2(new_n684_), .A3(new_n544_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G36gat), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n525_), .A2(G36gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n555_), .A2(new_n665_), .A3(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT45), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n689_), .A2(KEYINPUT46), .A3(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1329gat));
  NAND4_X1  g496(.A1(new_n680_), .A2(new_n684_), .A3(G43gat), .A4(new_n541_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n666_), .A2(new_n548_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(G43gat), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g500(.A(G50gat), .B1(new_n667_), .B2(new_n543_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n543_), .A2(G50gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n685_), .B2(new_n703_), .ZN(G1331gat));
  INV_X1    g503(.A(new_n279_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n315_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(new_n554_), .A3(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n631_), .ZN(new_n708_));
  INV_X1    g507(.A(G57gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n476_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n279_), .A2(new_n571_), .A3(new_n319_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n637_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G57gat), .B1(new_n712_), .B2(new_n527_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(G1332gat));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n708_), .A2(new_n715_), .A3(new_n544_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n712_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n544_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(G64gat), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G64gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT111), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n724_), .B(new_n716_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1333gat));
  INV_X1    g525(.A(G71gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n708_), .A2(new_n727_), .A3(new_n541_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT49), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n717_), .A2(new_n541_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(G71gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT49), .B(new_n727_), .C1(new_n717_), .C2(new_n541_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT112), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n735_), .B(new_n728_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1334gat));
  OAI21_X1  g536(.A(G78gat), .B1(new_n712_), .B2(new_n518_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT50), .ZN(new_n739_));
  INV_X1    g538(.A(G78gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n708_), .A2(new_n740_), .A3(new_n543_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1335gat));
  NOR2_X1   g541(.A1(new_n315_), .A2(new_n570_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n678_), .A2(new_n705_), .A3(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G85gat), .B1(new_n744_), .B2(new_n527_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n707_), .A2(new_n665_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n220_), .A3(new_n476_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1336gat));
  OAI21_X1  g547(.A(G92gat), .B1(new_n744_), .B2(new_n525_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n746_), .A2(new_n221_), .A3(new_n544_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1337gat));
  OAI21_X1  g550(.A(G99gat), .B1(new_n744_), .B2(new_n548_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n746_), .A2(new_n210_), .A3(new_n211_), .A4(new_n541_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g554(.A1(new_n746_), .A2(new_n209_), .A3(new_n543_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n705_), .A2(new_n743_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n682_), .A2(new_n757_), .ZN(new_n758_));
  AOI211_X1 g557(.A(KEYINPUT52), .B(new_n234_), .C1(new_n758_), .C2(new_n543_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n678_), .A2(new_n543_), .A3(new_n705_), .A4(new_n743_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(G106gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n756_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n756_), .C1(new_n759_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  NOR3_X1   g566(.A1(new_n319_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n570_), .B(new_n768_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n769_), .A2(KEYINPUT115), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n631_), .A2(KEYINPUT114), .A3(new_n768_), .A4(new_n770_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n293_), .A2(new_n294_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT119), .B1(new_n781_), .B2(new_n307_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n294_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n299_), .B2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(KEYINPUT119), .A3(new_n307_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n308_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n273_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n256_), .A2(new_n259_), .A3(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n258_), .A2(new_n252_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n255_), .B(new_n247_), .C1(new_n245_), .C2(KEYINPUT12), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n790_), .A2(KEYINPUT55), .B1(new_n250_), .B2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n272_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n793_), .A2(KEYINPUT56), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(KEYINPUT56), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n787_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT58), .B1(new_n796_), .B2(KEYINPUT120), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT120), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n793_), .B(KEYINPUT56), .Z(new_n800_));
  OAI211_X1 g599(.A(new_n798_), .B(new_n799_), .C1(new_n800_), .C2(new_n787_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n626_), .A2(new_n630_), .A3(new_n797_), .A4(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n271_), .A2(new_n273_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(new_n786_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n795_), .A2(KEYINPUT118), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n793_), .A2(new_n807_), .A3(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n793_), .A2(KEYINPUT116), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n793_), .B2(KEYINPUT116), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n806_), .B(new_n808_), .C1(new_n810_), .C2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n315_), .A2(new_n273_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n805_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n636_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n803_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n808_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n807_), .B1(new_n793_), .B2(KEYINPUT56), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n793_), .A2(KEYINPUT116), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n814_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT57), .B(new_n636_), .C1(new_n824_), .C2(new_n805_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n802_), .A2(new_n818_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n570_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n802_), .A2(new_n818_), .A3(KEYINPUT121), .A4(new_n825_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n776_), .A2(new_n780_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n545_), .A2(new_n541_), .A3(new_n476_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(G113gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n315_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT59), .B1(new_n830_), .B2(new_n831_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n831_), .A2(KEYINPUT59), .ZN(new_n836_));
  INV_X1    g635(.A(new_n825_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n802_), .A2(new_n818_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n802_), .A2(new_n818_), .A3(KEYINPUT122), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n570_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n774_), .A2(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n836_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n835_), .A2(new_n319_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n834_), .B1(new_n846_), .B2(new_n833_), .ZN(G1340gat));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n844_), .A2(new_n705_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n826_), .A2(new_n827_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n571_), .A3(new_n829_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n780_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n769_), .A2(KEYINPUT115), .A3(new_n771_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT115), .B1(new_n769_), .B2(new_n771_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n852_), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n831_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n850_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n848_), .B1(new_n849_), .B2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n835_), .A2(KEYINPUT123), .A3(new_n705_), .A4(new_n844_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(G120gat), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n279_), .B2(KEYINPUT60), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n832_), .B(new_n864_), .C1(KEYINPUT60), .C2(new_n863_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1341gat));
  INV_X1    g665(.A(G127gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n832_), .A2(new_n867_), .A3(new_n570_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n835_), .A2(new_n570_), .A3(new_n844_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n870_), .B2(new_n867_), .ZN(G1342gat));
  INV_X1    g670(.A(G134gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n832_), .A2(new_n872_), .A3(new_n817_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n669_), .A2(new_n670_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n835_), .A2(new_n874_), .A3(new_n844_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n873_), .B1(new_n876_), .B2(new_n872_), .ZN(G1343gat));
  NAND3_X1  g676(.A1(new_n526_), .A2(new_n548_), .A3(new_n476_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT124), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n857_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n315_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n705_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT125), .B(G148gat), .Z(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1345gat));
  NAND3_X1  g684(.A1(new_n857_), .A2(new_n570_), .A3(new_n879_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT126), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n857_), .A2(new_n888_), .A3(new_n570_), .A4(new_n879_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT61), .B(G155gat), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n887_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1346gat));
  AOI21_X1  g692(.A(G162gat), .B1(new_n880_), .B2(new_n817_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n671_), .A2(new_n673_), .A3(G162gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n880_), .B2(new_n895_), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n525_), .A2(new_n476_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n548_), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n518_), .B(new_n899_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900_), .B2(new_n706_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n842_), .A2(new_n843_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n543_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n905_), .A2(new_n385_), .A3(new_n315_), .A4(new_n899_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT62), .B(G169gat), .C1(new_n900_), .C2(new_n706_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n903_), .A2(new_n906_), .A3(new_n907_), .ZN(G1348gat));
  OR2_X1    g707(.A1(new_n900_), .A2(new_n279_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n830_), .A2(new_n543_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n899_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n279_), .A2(new_n386_), .A3(new_n911_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n909_), .A2(new_n386_), .B1(new_n910_), .B2(new_n912_), .ZN(G1349gat));
  NAND3_X1  g712(.A1(new_n910_), .A2(new_n570_), .A3(new_n899_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n911_), .A2(new_n571_), .A3(new_n401_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n914_), .A2(new_n420_), .B1(new_n905_), .B2(new_n915_), .ZN(G1350gat));
  INV_X1    g715(.A(new_n874_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G190gat), .B1(new_n900_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n817_), .A2(new_n400_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n900_), .B2(new_n919_), .ZN(G1351gat));
  NOR3_X1   g719(.A1(new_n898_), .A2(new_n541_), .A3(new_n518_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n857_), .A2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n315_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g724(.A1(new_n922_), .A2(new_n279_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT127), .B(G204gat), .Z(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n926_), .B2(new_n929_), .ZN(G1353gat));
  AOI211_X1 g729(.A(KEYINPUT63), .B(G211gat), .C1(new_n923_), .C2(new_n570_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT63), .B(G211gat), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n922_), .A2(new_n571_), .A3(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1354gat));
  OR3_X1    g733(.A1(new_n922_), .A2(G218gat), .A3(new_n636_), .ZN(new_n935_));
  OAI21_X1  g734(.A(G218gat), .B1(new_n922_), .B2(new_n917_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1355gat));
endmodule


