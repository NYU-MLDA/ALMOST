//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_;
  INV_X1    g000(.A(KEYINPUT24), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT82), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT82), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(G169gat), .B2(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT83), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n202_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n205_), .A2(new_n207_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT83), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n202_), .B1(G169gat), .B2(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT23), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT84), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT25), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n225_), .A2(KEYINPUT25), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228_));
  OR2_X1    g027(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n226_), .B(new_n227_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n211_), .A2(new_n216_), .A3(new_n224_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n203_), .A2(KEYINPUT22), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT22), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G169gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n237_), .A3(new_n204_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n229_), .A2(new_n225_), .A3(new_n230_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n218_), .A2(new_n223_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n234_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT30), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G71gat), .B(G99gat), .ZN(new_n247_));
  INV_X1    g046(.A(G43gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G15gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n249_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n246_), .B(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT85), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G127gat), .B(G134gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT31), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n254_), .B(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT2), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT2), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT3), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n262_), .A2(new_n264_), .A3(new_n265_), .A4(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G155gat), .ZN(new_n270_));
  INV_X1    g069(.A(G162gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(KEYINPUT86), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(G155gat), .B2(G162gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT87), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT87), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(G155gat), .A3(G162gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n269_), .A2(new_n275_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n275_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT88), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT88), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n277_), .A2(new_n279_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n275_), .B(new_n287_), .C1(new_n288_), .C2(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n284_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n261_), .A2(new_n266_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n282_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT97), .ZN(new_n294_));
  INV_X1    g093(.A(new_n257_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n294_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n257_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n296_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G225gat), .A2(G233gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT4), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n291_), .A2(new_n292_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n281_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT97), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(new_n297_), .A3(new_n257_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n303_), .B1(new_n307_), .B2(new_n296_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n301_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n257_), .A2(KEYINPUT4), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n293_), .B2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n302_), .B1(new_n308_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G29gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT0), .ZN(new_n315_));
  INV_X1    g114(.A(G57gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G85gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n302_), .B(new_n318_), .C1(new_n308_), .C2(new_n312_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n259_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n324_), .B1(new_n293_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT93), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n293_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G78gat), .B(G106gat), .ZN(new_n333_));
  INV_X1    g132(.A(G228gat), .ZN(new_n334_));
  INV_X1    g133(.A(G233gat), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n335_), .A2(KEYINPUT89), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(KEYINPUT89), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT90), .ZN(new_n339_));
  INV_X1    g138(.A(new_n292_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n280_), .A2(KEYINPUT1), .B1(new_n274_), .B2(new_n272_), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n341_), .A2(new_n287_), .B1(new_n284_), .B2(new_n288_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n340_), .B1(new_n342_), .B2(new_n286_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT29), .B1(new_n343_), .B2(new_n282_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT21), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n345_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(G197gat), .A2(G204gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(KEYINPUT21), .A3(new_n346_), .ZN(new_n351_));
  INV_X1    g150(.A(G211gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G218gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT91), .ZN(new_n354_));
  INV_X1    g153(.A(G218gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(G211gat), .B2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n349_), .A2(new_n351_), .A3(new_n353_), .A4(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(G211gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n353_), .A2(new_n358_), .A3(KEYINPUT91), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n359_), .A2(KEYINPUT21), .A3(new_n350_), .A4(new_n346_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n339_), .B1(new_n344_), .B2(new_n361_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n357_), .A2(new_n360_), .A3(KEYINPUT92), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT92), .B1(new_n357_), .B2(new_n360_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n339_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(KEYINPUT29), .B2(new_n305_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n333_), .B1(new_n362_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n361_), .B1(new_n293_), .B2(new_n325_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n339_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n344_), .A2(new_n339_), .A3(new_n365_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n333_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G22gat), .B(G50gat), .Z(new_n375_));
  AND3_X1   g174(.A1(new_n368_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n332_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n375_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n362_), .A2(new_n367_), .A3(new_n333_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n373_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n368_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n330_), .A2(new_n331_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT20), .B1(new_n245_), .B2(new_n365_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n361_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT95), .ZN(new_n392_));
  INV_X1    g191(.A(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n225_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n239_), .B1(new_n224_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n212_), .A2(new_n202_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT26), .B(G190gat), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n396_), .A2(new_n398_), .A3(new_n242_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n392_), .A2(new_n395_), .B1(new_n399_), .B2(new_n216_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n224_), .A2(new_n394_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n240_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT95), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n391_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n389_), .B1(new_n390_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n245_), .A2(new_n365_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n389_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n407_), .A2(KEYINPUT20), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n400_), .A2(new_n403_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n406_), .B(new_n408_), .C1(new_n409_), .C2(new_n361_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n405_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G8gat), .B(G36gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(G64gat), .B(G92gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n405_), .A2(new_n410_), .A3(new_n416_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT27), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(KEYINPUT27), .ZN(new_n421_));
  INV_X1    g220(.A(new_n390_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n409_), .A2(new_n361_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n407_), .A3(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT99), .B(KEYINPUT20), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n395_), .A2(new_n361_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n399_), .A2(new_n216_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n407_), .B1(new_n406_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n416_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT102), .B1(new_n421_), .B2(new_n431_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n390_), .A2(new_n404_), .A3(new_n389_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n417_), .B1(new_n433_), .B2(new_n429_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT102), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(KEYINPUT27), .A4(new_n419_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n420_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT103), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n386_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n386_), .B2(new_n437_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n323_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT104), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT104), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(new_n323_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT101), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n320_), .A2(new_n321_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n416_), .A2(KEYINPUT32), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n405_), .A2(new_n410_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n424_), .A2(new_n430_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n447_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n449_), .A2(KEYINPUT100), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT100), .B1(new_n449_), .B2(new_n450_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n448_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n445_), .B1(new_n446_), .B2(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n451_), .A2(new_n452_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n455_), .A2(new_n322_), .A3(KEYINPUT101), .A4(new_n448_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n418_), .A2(new_n419_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n308_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n458_), .B(new_n301_), .C1(new_n293_), .C2(new_n311_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n318_), .B1(new_n300_), .B2(new_n309_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n457_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT98), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n321_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT33), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n321_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n454_), .A2(new_n456_), .A3(new_n467_), .A4(new_n386_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n259_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n446_), .A2(new_n437_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n386_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n442_), .A2(new_n444_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT13), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT71), .ZN(new_n476_));
  OR2_X1    g275(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(G78gat), .ZN(new_n480_));
  INV_X1    g279(.A(G78gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(new_n481_), .A3(new_n478_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G57gat), .B(G64gat), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n480_), .A2(new_n482_), .B1(KEYINPUT11), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n482_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n483_), .B(KEYINPUT11), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n484_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G85gat), .B(G92gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(G99gat), .ZN(new_n491_));
  INV_X1    g290(.A(G106gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(KEYINPUT7), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(G99gat), .B2(G106gat), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n490_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT67), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT8), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT65), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n493_), .A2(new_n495_), .ZN(new_n506_));
  AND3_X1   g305(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n506_), .A2(new_n509_), .A3(KEYINPUT65), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT66), .B(KEYINPUT8), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n489_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n505_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n489_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT67), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n503_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  AND2_X1   g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(KEYINPUT9), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT64), .B(G85gat), .Z(new_n521_));
  INV_X1    g320(.A(G92gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n520_), .B1(new_n523_), .B2(KEYINPUT9), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT10), .B(G99gat), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n524_), .B(new_n509_), .C1(G106gat), .C2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n488_), .B1(new_n517_), .B2(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n527_), .A2(KEYINPUT69), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n517_), .A2(new_n526_), .A3(new_n488_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(new_n527_), .B2(KEYINPUT69), .ZN(new_n530_));
  OAI211_X1 g329(.A(G230gat), .B(G233gat), .C1(new_n528_), .C2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n517_), .A2(new_n526_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n488_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT12), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT70), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n535_), .A2(KEYINPUT70), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n536_), .B1(new_n527_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G230gat), .A2(G233gat), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n538_), .A2(new_n540_), .A3(new_n541_), .A4(new_n529_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n531_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G120gat), .B(G148gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT5), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G176gat), .B(G204gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  OAI21_X1  g346(.A(new_n476_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n531_), .A2(KEYINPUT71), .A3(new_n542_), .A4(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n543_), .A2(new_n547_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n551_), .A2(KEYINPUT72), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT72), .B1(new_n551_), .B2(new_n552_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n475_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n552_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n551_), .A2(KEYINPUT72), .A3(new_n552_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(KEYINPUT13), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G29gat), .B(G36gat), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT73), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G43gat), .B(G50gat), .Z(new_n566_));
  OR3_X1    g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT80), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT77), .B(G1gat), .ZN(new_n571_));
  INV_X1    g370(.A(G8gat), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT14), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G15gat), .B(G22gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G1gat), .B(G8gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n570_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n577_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n570_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT15), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n569_), .B(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n577_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n579_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n581_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G113gat), .B(G141gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G169gat), .B(G197gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n581_), .A2(new_n588_), .A3(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n561_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n474_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT74), .ZN(new_n601_));
  XOR2_X1   g400(.A(G134gat), .B(G162gat), .Z(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n585_), .A2(new_n532_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n532_), .A2(new_n569_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT34), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT35), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n607_), .A2(new_n608_), .A3(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n611_), .A2(new_n612_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n607_), .A2(new_n617_), .A3(new_n608_), .A4(new_n613_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT75), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n606_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n616_), .A2(KEYINPUT75), .A3(new_n605_), .A4(new_n618_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n603_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(KEYINPUT36), .A3(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n621_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT76), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(KEYINPUT37), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n621_), .A2(new_n624_), .A3(new_n622_), .A4(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n488_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(new_n582_), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT79), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G127gat), .B(G155gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G183gat), .B(G211gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n636_), .B(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT17), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n640_), .A2(new_n641_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n634_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n634_), .A2(new_n642_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n631_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n599_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n571_), .A3(new_n322_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT105), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n555_), .A2(new_n560_), .A3(new_n646_), .A4(new_n596_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n625_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n474_), .A2(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n322_), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n650_), .A2(new_n651_), .B1(new_n660_), .B2(G1gat), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n653_), .A2(new_n661_), .ZN(G1324gat));
  INV_X1    g461(.A(new_n437_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n649_), .A2(new_n572_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n656_), .A2(new_n658_), .A3(new_n663_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(G8gat), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n666_), .A2(new_n665_), .A3(G8gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n664_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT40), .B(new_n664_), .C1(new_n669_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1325gat));
  NAND2_X1  g475(.A1(new_n659_), .A2(new_n469_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G15gat), .ZN(new_n678_));
  XOR2_X1   g477(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n679_));
  OR2_X1    g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n679_), .ZN(new_n681_));
  INV_X1    g480(.A(G15gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n649_), .A2(new_n682_), .A3(new_n469_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n681_), .A3(new_n683_), .ZN(G1326gat));
  INV_X1    g483(.A(G22gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n649_), .A2(new_n685_), .A3(new_n471_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n659_), .A2(new_n471_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(G22gat), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT42), .B(new_n685_), .C1(new_n659_), .C2(new_n471_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT109), .ZN(G1327gat));
  NOR2_X1   g491(.A1(new_n657_), .A2(new_n646_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n599_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n322_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n598_), .A2(new_n647_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n631_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n698_), .B2(KEYINPUT110), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n474_), .B2(new_n631_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n474_), .A2(new_n631_), .A3(new_n699_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n697_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT44), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n704_), .A2(G29gat), .A3(new_n322_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n703_), .A2(KEYINPUT44), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n696_), .B1(new_n705_), .B2(new_n706_), .ZN(G1328gat));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n695_), .A2(new_n708_), .A3(new_n663_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT45), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n437_), .B1(new_n703_), .B2(KEYINPUT44), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n706_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n710_), .B(KEYINPUT46), .C1(new_n712_), .C2(new_n708_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n709_), .B(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n708_), .B1(new_n706_), .B2(new_n711_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n714_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n713_), .A2(new_n718_), .ZN(G1329gat));
  OAI21_X1  g518(.A(new_n248_), .B1(new_n694_), .B2(new_n259_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n704_), .A2(G43gat), .A3(new_n469_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n703_), .A2(KEYINPUT44), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n695_), .B2(new_n471_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n704_), .A2(G50gat), .A3(new_n471_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n706_), .ZN(G1331gat));
  NAND2_X1  g526(.A1(new_n561_), .A2(new_n648_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT111), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n474_), .A2(new_n597_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n316_), .B1(new_n731_), .B2(new_n446_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n733_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n596_), .A2(new_n647_), .ZN(new_n736_));
  AND4_X1   g535(.A1(new_n657_), .A2(new_n474_), .A3(new_n561_), .A4(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(G57gat), .A3(new_n322_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n734_), .A2(new_n735_), .A3(new_n738_), .ZN(G1332gat));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n663_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G64gat), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n742_));
  OR2_X1    g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n742_), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n731_), .A2(G64gat), .A3(new_n437_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n737_), .B2(new_n469_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT49), .Z(new_n749_));
  NAND2_X1  g548(.A1(new_n469_), .A2(new_n747_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT114), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n731_), .B2(new_n751_), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n737_), .A2(new_n471_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G78gat), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(KEYINPUT50), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(KEYINPUT50), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n471_), .A2(new_n481_), .ZN(new_n757_));
  OAI22_X1  g556(.A1(new_n755_), .A2(new_n756_), .B1(new_n731_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT115), .ZN(G1335gat));
  AND3_X1   g558(.A1(new_n730_), .A2(new_n561_), .A3(new_n693_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n322_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n701_), .A2(new_n702_), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n646_), .B(new_n596_), .C1(new_n555_), .C2(new_n560_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n446_), .A2(new_n521_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n761_), .B1(new_n765_), .B2(new_n766_), .ZN(G1336gat));
  OAI21_X1  g566(.A(G92gat), .B1(new_n764_), .B2(new_n437_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n760_), .A2(new_n522_), .A3(new_n663_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1337gat));
  NOR2_X1   g569(.A1(new_n259_), .A2(new_n525_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n760_), .A2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT116), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n491_), .B1(new_n765_), .B2(new_n469_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT51), .B1(new_n773_), .B2(new_n776_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1338gat));
  AND3_X1   g579(.A1(new_n474_), .A2(new_n631_), .A3(new_n699_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n471_), .B(new_n763_), .C1(new_n781_), .C2(new_n700_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(G106gat), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT117), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n782_), .A2(new_n786_), .A3(new_n783_), .A4(G106gat), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n782_), .A2(G106gat), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT52), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n785_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n760_), .A2(new_n492_), .A3(new_n471_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT53), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n790_), .A2(new_n794_), .A3(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n583_), .A2(new_n586_), .A3(new_n580_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n592_), .B(new_n797_), .C1(new_n578_), .C2(new_n580_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n594_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n542_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n529_), .B1(new_n527_), .B2(new_n536_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n804_), .A2(KEYINPUT55), .A3(new_n541_), .A4(new_n540_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n539_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n537_), .B1(new_n534_), .B2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(G230gat), .B(G233gat), .C1(new_n807_), .C2(new_n803_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n802_), .A2(new_n805_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT119), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n802_), .A2(new_n805_), .A3(new_n811_), .A4(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n547_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n815_), .B(new_n549_), .C1(new_n810_), .C2(new_n812_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n800_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT58), .B(new_n800_), .C1(new_n814_), .C2(new_n816_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n631_), .A3(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n596_), .A2(new_n551_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n799_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n625_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n821_), .B1(KEYINPUT57), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(KEYINPUT57), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n647_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n627_), .A2(new_n630_), .A3(new_n736_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n560_), .A3(new_n555_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT54), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT118), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n832_), .A2(new_n835_), .A3(KEYINPUT54), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n834_), .B(new_n836_), .C1(KEYINPUT54), .C2(new_n832_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n830_), .A2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n322_), .B(new_n469_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT59), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n832_), .A2(KEYINPUT54), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n834_), .A2(new_n836_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n549_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT56), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT58), .B1(new_n847_), .B2(new_n800_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n820_), .A2(new_n631_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n823_), .A2(new_n825_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT57), .B1(new_n851_), .B2(new_n657_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n845_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n821_), .B(KEYINPUT120), .C1(KEYINPUT57), .C2(new_n826_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n828_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n844_), .B1(new_n855_), .B2(new_n647_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n839_), .A2(KEYINPUT59), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n842_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n597_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n597_), .A2(G113gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n841_), .B2(new_n860_), .ZN(G1340gat));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n862_));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n561_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n838_), .A2(new_n840_), .A3(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n842_), .B(new_n561_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n866_), .B1(new_n868_), .B2(new_n863_), .ZN(G1341gat));
  OAI21_X1  g668(.A(G127gat), .B1(new_n858_), .B2(new_n647_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n647_), .A2(G127gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n841_), .B2(new_n871_), .ZN(G1342gat));
  OAI21_X1  g671(.A(G134gat), .B1(new_n858_), .B2(new_n698_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n657_), .A2(G134gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n841_), .B2(new_n874_), .ZN(G1343gat));
  INV_X1    g674(.A(new_n838_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n469_), .A2(new_n386_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n437_), .A3(new_n322_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n596_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n561_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n646_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  NOR2_X1   g685(.A1(new_n657_), .A2(G162gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n879_), .A2(new_n887_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n876_), .A2(new_n698_), .A3(new_n878_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n271_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT121), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n888_), .B(new_n892_), .C1(new_n271_), .C2(new_n889_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1347gat));
  NOR3_X1   g693(.A1(new_n259_), .A2(new_n437_), .A3(new_n322_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n856_), .A2(new_n471_), .A3(new_n896_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n897_), .A2(new_n596_), .A3(new_n235_), .A4(new_n237_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n596_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT122), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n900_), .A2(KEYINPUT122), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n902_), .A2(new_n903_), .A3(new_n471_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n855_), .A2(new_n647_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n837_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n203_), .B1(new_n907_), .B2(KEYINPUT123), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n856_), .B2(new_n905_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n899_), .B1(new_n908_), .B2(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n829_), .B1(new_n827_), .B2(new_n845_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n646_), .B1(new_n912_), .B2(new_n854_), .ZN(new_n913_));
  OAI211_X1 g712(.A(KEYINPUT123), .B(new_n904_), .C1(new_n913_), .C2(new_n844_), .ZN(new_n914_));
  AND4_X1   g713(.A1(new_n899_), .A2(new_n910_), .A3(new_n914_), .A4(G169gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n898_), .B1(new_n911_), .B2(new_n915_), .ZN(G1348gat));
  NAND3_X1  g715(.A1(new_n561_), .A2(G176gat), .A3(new_n895_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n876_), .A2(new_n471_), .A3(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n896_), .A2(new_n471_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n561_), .B(new_n919_), .C1(new_n913_), .C2(new_n844_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n204_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n920_), .A2(KEYINPUT124), .A3(new_n204_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n918_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  NAND2_X1  g724(.A1(new_n227_), .A2(new_n226_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n646_), .A2(new_n926_), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n856_), .A2(new_n471_), .A3(new_n896_), .A4(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n896_), .A2(new_n647_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n838_), .A2(new_n386_), .A3(new_n929_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n930_), .A2(new_n225_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n928_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT125), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n934_), .B1(new_n928_), .B2(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n897_), .A2(new_n625_), .A3(new_n397_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n897_), .A2(new_n631_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n393_), .ZN(G1351gat));
  NOR3_X1   g738(.A1(new_n469_), .A2(new_n386_), .A3(new_n322_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n940_), .A2(KEYINPUT126), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(KEYINPUT126), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n941_), .A2(new_n942_), .A3(new_n437_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n838_), .A2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n596_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n561_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g748(.A1(new_n944_), .A2(new_n647_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  AND2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n950_), .B1(new_n951_), .B2(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n953_), .B1(new_n950_), .B2(new_n951_), .ZN(G1354gat));
  OAI21_X1  g753(.A(G218gat), .B1(new_n944_), .B2(new_n698_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n625_), .A2(new_n355_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n944_), .B2(new_n956_), .ZN(G1355gat));
endmodule


