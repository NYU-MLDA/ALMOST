//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G230gat), .A2(G233gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208_));
  INV_X1    g007(.A(G57gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G64gat), .ZN(new_n210_));
  INV_X1    g009(.A(G64gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(G57gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n208_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(G57gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n209_), .A2(G64gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT66), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G71gat), .B(G78gat), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n213_), .A2(new_n217_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(KEYINPUT11), .ZN(new_n223_));
  AOI211_X1 g022(.A(KEYINPUT67), .B(new_n214_), .C1(new_n213_), .C2(new_n217_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n220_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  INV_X1    g027(.A(G106gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT6), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(KEYINPUT6), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n226_), .B(new_n230_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  XOR2_X1   g035(.A(G85gat), .B(G92gat), .Z(new_n237_));
  AND3_X1   g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n236_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT65), .B(G92gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT64), .B(G85gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT9), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G85gat), .ZN(new_n244_));
  INV_X1    g043(.A(G92gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT9), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n243_), .A2(new_n246_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT10), .B(G99gat), .Z(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n229_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n249_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n250_));
  OAI22_X1  g049(.A1(new_n238_), .A2(new_n239_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT66), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(new_n215_), .B2(new_n216_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT11), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT67), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n222_), .A2(new_n221_), .A3(KEYINPUT11), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n225_), .A2(new_n251_), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n251_), .B1(new_n257_), .B2(new_n225_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n207_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(KEYINPUT68), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(KEYINPUT68), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT12), .B1(new_n258_), .B2(new_n259_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n225_), .A2(new_n251_), .A3(new_n257_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n206_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n205_), .B1(new_n263_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n205_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n261_), .A2(new_n268_), .A3(new_n262_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT13), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(KEYINPUT13), .A3(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G113gat), .B(G141gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT79), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G169gat), .B(G197gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G229gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT75), .ZN(new_n284_));
  INV_X1    g083(.A(G22gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(KEYINPUT71), .A2(G15gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(KEYINPUT71), .A2(G15gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n285_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n290_));
  INV_X1    g089(.A(G15gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(G22gat), .A3(new_n286_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT14), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n295_), .B1(G1gat), .B2(G8gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G8gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n294_), .A2(new_n301_), .A3(new_n297_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G29gat), .B(G36gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G43gat), .B(G50gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n284_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n310_));
  AOI211_X1 g109(.A(KEYINPUT76), .B(new_n306_), .C1(new_n300_), .C2(new_n302_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n308_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n301_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n313_));
  AOI211_X1 g112(.A(new_n296_), .B(new_n299_), .C1(new_n289_), .C2(new_n293_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT75), .B1(new_n315_), .B2(new_n306_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT76), .B1(new_n315_), .B2(new_n306_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n303_), .A2(new_n309_), .A3(new_n307_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n283_), .B1(new_n312_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n307_), .A2(KEYINPUT15), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT15), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n306_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n303_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n315_), .A2(new_n306_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n283_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT77), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n320_), .A2(new_n328_), .ZN(new_n329_));
  AOI211_X1 g128(.A(KEYINPUT77), .B(new_n283_), .C1(new_n312_), .C2(new_n319_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n282_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(KEYINPUT80), .B(new_n282_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT78), .B1(new_n329_), .B2(new_n330_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n320_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n338_), .B(new_n339_), .C1(new_n320_), .C2(new_n328_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n340_), .A3(new_n281_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n342_), .A2(KEYINPUT81), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(KEYINPUT81), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT82), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(KEYINPUT24), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT83), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n350_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n347_), .A2(KEYINPUT24), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT25), .B(G183gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(G190gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT23), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .A4(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G169gat), .ZN(new_n361_));
  INV_X1    g160(.A(G176gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n363_), .B(KEYINPUT84), .Z(new_n364_));
  OAI21_X1  g163(.A(new_n358_), .B1(G183gat), .B2(G190gat), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n365_), .A2(new_n348_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n360_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n360_), .A2(KEYINPUT85), .A3(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  INV_X1    g172(.A(G71gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(new_n228_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n372_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G15gat), .B(G43gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT86), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT30), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G127gat), .B(G134gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G113gat), .B(G120gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n382_), .B(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n379_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n366_), .A2(new_n363_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G211gat), .B(G218gat), .ZN(new_n393_));
  INV_X1    g192(.A(G197gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(G204gat), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n393_), .B(KEYINPUT21), .C1(KEYINPUT90), .C2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G197gat), .B(G204gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n393_), .A2(KEYINPUT21), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(new_n397_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n396_), .B2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n403_));
  NAND3_X1  g202(.A1(new_n347_), .A2(new_n348_), .A3(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n359_), .B(new_n404_), .C1(new_n347_), .C2(new_n403_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n392_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n406_));
  AOI211_X1 g205(.A(new_n389_), .B(new_n391_), .C1(new_n406_), .C2(KEYINPUT93), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n406_), .A2(KEYINPUT93), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n402_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n370_), .A2(new_n371_), .A3(new_n402_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n392_), .A2(new_n405_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n402_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n389_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n391_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT18), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  NAND3_X1  g220(.A1(new_n411_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n409_), .A2(new_n410_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n391_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n423_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT27), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n422_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT96), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n422_), .A2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n411_), .A2(new_n417_), .A3(KEYINPUT96), .A4(new_n421_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n406_), .A2(KEYINPUT20), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n391_), .B1(new_n410_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n391_), .B2(new_n416_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n423_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n431_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n429_), .B1(new_n437_), .B2(KEYINPUT27), .ZN(new_n438_));
  NOR2_X1   g237(.A1(G141gat), .A2(G148gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT3), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT2), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT89), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446_));
  OR2_X1    g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n439_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(KEYINPUT1), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n447_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n446_), .A2(KEYINPUT1), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n441_), .B(new_n449_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n453_), .B(KEYINPUT88), .Z(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n385_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT94), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n455_), .A2(KEYINPUT94), .A3(new_n456_), .A4(new_n385_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G225gat), .A2(G233gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n455_), .A2(new_n385_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n385_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n448_), .A2(new_n465_), .A3(new_n454_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(KEYINPUT4), .A3(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n464_), .A2(new_n466_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n462_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G1gat), .B(G29gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(G85gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT0), .B(G57gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(new_n474_), .Z(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n468_), .A2(new_n475_), .A3(new_n470_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(G50gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT28), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n455_), .B2(KEYINPUT29), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT29), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n448_), .A2(KEYINPUT28), .A3(new_n483_), .A4(new_n454_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n285_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n285_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n480_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G78gat), .B(G106gat), .ZN(new_n489_));
  INV_X1    g288(.A(G228gat), .ZN(new_n490_));
  INV_X1    g289(.A(G233gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n455_), .A2(KEYINPUT29), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n494_), .B2(new_n414_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n483_), .B1(new_n448_), .B2(new_n454_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n496_), .A2(new_n492_), .A3(new_n402_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n489_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT91), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n482_), .A2(new_n484_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G22gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(G50gat), .A3(new_n485_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n488_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n489_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n497_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n492_), .B1(new_n496_), .B2(new_n402_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n495_), .A2(new_n497_), .A3(new_n489_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n507_), .A2(new_n508_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n511_), .A2(new_n499_), .A3(new_n502_), .A4(new_n488_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n438_), .A2(new_n479_), .A3(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n510_), .A2(new_n512_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n464_), .A2(new_n466_), .A3(new_n463_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n476_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n461_), .A2(new_n467_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n518_), .B2(new_n462_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT33), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n478_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n478_), .A2(new_n520_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n422_), .A4(new_n427_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n421_), .A2(KEYINPUT32), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT95), .B1(new_n435_), .B2(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n424_), .A2(new_n426_), .A3(new_n525_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n435_), .A2(KEYINPUT95), .A3(new_n525_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n479_), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n515_), .B1(new_n523_), .B2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n388_), .B1(new_n514_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT97), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n438_), .B2(new_n515_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n479_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n422_), .A2(new_n430_), .B1(new_n435_), .B2(new_n423_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n428_), .B1(new_n536_), .B2(new_n432_), .ZN(new_n537_));
  OAI211_X1 g336(.A(KEYINPUT97), .B(new_n513_), .C1(new_n537_), .C2(new_n429_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n534_), .A2(new_n535_), .A3(new_n387_), .A4(new_n538_), .ZN(new_n539_));
  AOI211_X1 g338(.A(new_n277_), .B(new_n345_), .C1(new_n532_), .C2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n247_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n250_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n233_), .B(new_n231_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n230_), .A2(new_n226_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n237_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT8), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n541_), .A2(new_n542_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n306_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n251_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT69), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n554_), .A2(new_n557_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n563_), .B(KEYINPUT36), .Z(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n565_), .A2(KEYINPUT37), .A3(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n560_), .A2(KEYINPUT70), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n560_), .A2(KEYINPUT70), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n566_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n565_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n568_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n315_), .B(new_n576_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n223_), .A2(new_n224_), .A3(new_n220_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n255_), .A2(new_n256_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n577_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT74), .B(KEYINPUT17), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n583_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT73), .B(KEYINPUT17), .Z(new_n590_));
  OR2_X1    g389(.A1(new_n581_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n575_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n540_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT98), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n540_), .A2(new_n597_), .A3(new_n594_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(G1gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n479_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT38), .ZN(new_n602_));
  INV_X1    g401(.A(new_n277_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n342_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT99), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(new_n593_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n571_), .A2(new_n565_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n532_), .B2(new_n539_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n535_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT100), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n602_), .A2(new_n611_), .ZN(G1324gat));
  INV_X1    g411(.A(new_n438_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(G8gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n596_), .A2(new_n598_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT101), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n596_), .A2(new_n617_), .A3(new_n598_), .A4(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  OAI221_X1 g420(.A(G8gat), .B1(new_n620_), .B2(new_n621_), .C1(new_n609_), .C2(new_n613_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n621_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n619_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n619_), .B2(new_n624_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(G1325gat));
  NAND3_X1  g427(.A1(new_n599_), .A2(new_n291_), .A3(new_n387_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n609_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n291_), .B1(new_n630_), .B2(new_n387_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n632_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n629_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT104), .ZN(G1326gat));
  NAND3_X1  g435(.A1(new_n599_), .A2(new_n285_), .A3(new_n515_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G22gat), .B1(new_n609_), .B2(new_n513_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1327gat));
  NOR2_X1   g439(.A1(new_n572_), .A2(new_n592_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n540_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n479_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n532_), .A2(new_n539_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n575_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT43), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n644_), .A2(new_n647_), .A3(new_n575_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n605_), .A2(new_n592_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n649_), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n647_), .B1(new_n644_), .B2(new_n575_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT43), .B(new_n574_), .C1(new_n532_), .C2(new_n539_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT44), .B(new_n650_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n649_), .A2(new_n650_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n651_), .A2(new_n656_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n479_), .A2(G29gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n643_), .B1(new_n659_), .B2(new_n660_), .ZN(G1328gat));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  INV_X1    g461(.A(G36gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n659_), .B2(new_n438_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n642_), .A2(new_n663_), .A3(new_n438_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT45), .Z(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n651_), .A2(new_n656_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n657_), .A2(new_n658_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n438_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G36gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n665_), .B(KEYINPUT45), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(KEYINPUT46), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n667_), .A2(new_n673_), .ZN(G1329gat));
  NAND4_X1  g473(.A1(new_n668_), .A2(G43gat), .A3(new_n387_), .A4(new_n669_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n642_), .A2(new_n387_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(G43gat), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n675_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1330gat));
  AOI21_X1  g482(.A(G50gat), .B1(new_n642_), .B2(new_n515_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n513_), .A2(new_n480_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n659_), .B2(new_n685_), .ZN(G1331gat));
  AOI211_X1 g485(.A(new_n342_), .B(new_n603_), .C1(new_n532_), .C2(new_n539_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(new_n594_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G57gat), .B1(new_n688_), .B2(new_n479_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT107), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n608_), .A2(new_n592_), .A3(new_n277_), .A4(new_n345_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n691_), .A2(new_n209_), .A3(new_n535_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT108), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n690_), .A2(new_n693_), .ZN(G1332gat));
  OAI21_X1  g493(.A(G64gat), .B1(new_n691_), .B2(new_n613_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT48), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n688_), .A2(new_n211_), .A3(new_n438_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1333gat));
  OAI21_X1  g497(.A(G71gat), .B1(new_n691_), .B2(new_n388_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT49), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n688_), .A2(new_n374_), .A3(new_n387_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1334gat));
  OAI21_X1  g501(.A(G78gat), .B1(new_n691_), .B2(new_n513_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT50), .ZN(new_n704_));
  INV_X1    g503(.A(G78gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n688_), .A2(new_n705_), .A3(new_n515_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1335gat));
  AND2_X1   g506(.A1(new_n687_), .A2(new_n641_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n479_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n244_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n710_), .A2(KEYINPUT109), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(KEYINPUT109), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n603_), .A2(new_n592_), .A3(new_n342_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n649_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(new_n479_), .A3(new_n241_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n711_), .A2(new_n712_), .A3(new_n715_), .ZN(G1336gat));
  AOI21_X1  g515(.A(G92gat), .B1(new_n708_), .B2(new_n438_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n438_), .A2(new_n240_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n714_), .B2(new_n718_), .ZN(G1337gat));
  AOI21_X1  g518(.A(new_n228_), .B1(new_n714_), .B2(new_n387_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n387_), .A2(new_n248_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n708_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n723_));
  MUX2_X1   g522(.A(KEYINPUT51), .B(new_n723_), .S(KEYINPUT111), .Z(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n725_), .B1(new_n722_), .B2(new_n723_), .ZN(G1338gat));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n649_), .A2(new_n727_), .A3(new_n515_), .A4(new_n713_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n515_), .B(new_n713_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT113), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n728_), .A2(new_n730_), .A3(G106gat), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n708_), .A2(new_n229_), .A3(new_n515_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT112), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n728_), .A2(new_n730_), .A3(KEYINPUT52), .A4(G106gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n733_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT53), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT53), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n733_), .A2(new_n735_), .A3(new_n739_), .A4(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1339gat));
  AND2_X1   g540(.A1(new_n534_), .A2(new_n387_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n479_), .A3(new_n538_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n272_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n335_), .B2(new_n341_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n264_), .A2(new_n267_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(new_n207_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n548_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n266_), .B1(new_n749_), .B2(new_n265_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n265_), .A2(new_n266_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT114), .B1(new_n752_), .B2(new_n206_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754_));
  NOR4_X1   g553(.A1(new_n750_), .A2(new_n751_), .A3(new_n754_), .A4(new_n207_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n748_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n207_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT55), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n752_), .A2(KEYINPUT114), .A3(new_n206_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n268_), .A2(new_n754_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n756_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT56), .B1(new_n762_), .B2(new_n205_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n764_), .B(new_n271_), .C1(new_n756_), .C2(new_n761_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n745_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n312_), .A2(new_n319_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n283_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n281_), .C1(new_n283_), .C2(new_n326_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n335_), .A2(new_n273_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n607_), .B1(new_n766_), .B2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT115), .B1(new_n772_), .B2(KEYINPUT57), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n758_), .B1(new_n760_), .B2(new_n759_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n205_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n764_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n762_), .A2(KEYINPUT56), .A3(new_n205_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n770_), .B1(new_n781_), .B2(new_n745_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n774_), .B(new_n775_), .C1(new_n782_), .C2(new_n607_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n773_), .A2(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n335_), .A2(new_n769_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n272_), .C1(new_n763_), .C2(new_n765_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n787_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n781_), .A2(new_n272_), .A3(new_n785_), .A4(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n575_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n772_), .A2(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n593_), .B1(new_n784_), .B2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n575_), .A2(new_n277_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n345_), .A2(new_n795_), .A3(new_n796_), .A4(new_n592_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n343_), .A2(new_n592_), .A3(new_n344_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n603_), .A2(new_n574_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT54), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n797_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n743_), .B1(new_n794_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G113gat), .B1(new_n803_), .B2(new_n342_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT117), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n803_), .B2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n773_), .A2(new_n783_), .A3(new_n791_), .A4(new_n792_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n801_), .B1(new_n809_), .B2(new_n593_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT118), .B(KEYINPUT59), .C1(new_n810_), .C2(new_n743_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n775_), .B1(new_n782_), .B2(new_n607_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n791_), .A2(new_n812_), .A3(new_n792_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n801_), .B1(new_n813_), .B2(new_n593_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n743_), .A2(KEYINPUT59), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT119), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n813_), .A2(new_n593_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n818_), .B(new_n815_), .C1(new_n819_), .C2(new_n801_), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n808_), .A2(new_n811_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(G113gat), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n345_), .A2(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT120), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n805_), .B1(new_n821_), .B2(new_n824_), .ZN(G1340gat));
  INV_X1    g624(.A(G120gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n821_), .B2(new_n277_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n803_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n603_), .B2(KEYINPUT60), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n826_), .A2(KEYINPUT60), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(KEYINPUT121), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(KEYINPUT121), .B2(new_n829_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n828_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT122), .B1(new_n827_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n835_));
  INV_X1    g634(.A(new_n833_), .ZN(new_n836_));
  AOI221_X4 g635(.A(new_n603_), .B1(new_n817_), .B2(new_n820_), .C1(new_n808_), .C2(new_n811_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n835_), .B(new_n836_), .C1(new_n837_), .C2(new_n826_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n838_), .ZN(G1341gat));
  INV_X1    g638(.A(G127gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n803_), .A2(new_n840_), .A3(new_n592_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n821_), .A2(new_n592_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n840_), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n803_), .A2(new_n844_), .A3(new_n607_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n821_), .A2(new_n575_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n844_), .ZN(G1343gat));
  NOR2_X1   g646(.A1(new_n810_), .A2(new_n387_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n438_), .A2(new_n535_), .A3(new_n513_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n342_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n277_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  OR3_X1    g655(.A1(new_n850_), .A2(new_n593_), .A3(new_n856_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n850_), .B2(new_n593_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1346gat));
  AOI21_X1  g661(.A(G162gat), .B1(new_n851_), .B2(new_n607_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n575_), .A2(G162gat), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n864_), .B(KEYINPUT125), .Z(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n851_), .B2(new_n865_), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n814_), .A2(new_n515_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n613_), .A2(new_n479_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n387_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n867_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n342_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(G169gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT127), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n875_), .A2(new_n876_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(KEYINPUT127), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n876_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n880_), .B(new_n881_), .C1(new_n873_), .C2(new_n874_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n873_), .A2(new_n361_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n879_), .A2(new_n882_), .A3(new_n883_), .ZN(G1348gat));
  INV_X1    g683(.A(new_n871_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G176gat), .B1(new_n885_), .B2(new_n277_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n810_), .A2(new_n515_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n869_), .A2(new_n362_), .A3(new_n603_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1349gat));
  NOR2_X1   g688(.A1(new_n869_), .A2(new_n593_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G183gat), .B1(new_n887_), .B2(new_n890_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n869_), .A2(new_n354_), .A3(new_n593_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n867_), .B2(new_n892_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n871_), .B2(new_n574_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n607_), .A2(new_n355_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n871_), .B2(new_n895_), .ZN(G1351gat));
  NOR3_X1   g695(.A1(new_n613_), .A2(new_n479_), .A3(new_n513_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n848_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n872_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n394_), .ZN(G1352gat));
  INV_X1    g699(.A(new_n898_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n277_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n592_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  AND2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n904_), .B2(new_n905_), .ZN(G1354gat));
  OR3_X1    g707(.A1(new_n898_), .A2(G218gat), .A3(new_n572_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G218gat), .B1(new_n898_), .B2(new_n574_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1355gat));
endmodule


