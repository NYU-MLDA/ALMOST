//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_;
  INV_X1    g000(.A(G230gat), .ZN(new_n202_));
  INV_X1    g001(.A(G233gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G71gat), .B(G78gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT11), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n208_));
  INV_X1    g007(.A(new_n206_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n207_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT10), .B(G99gat), .Z(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT6), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  INV_X1    g020(.A(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT9), .A3(new_n219_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .A4(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n219_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(KEYINPUT64), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT64), .B1(new_n227_), .B2(KEYINPUT65), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT6), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n217_), .B(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(G99gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n215_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n229_), .B(new_n230_), .C1(new_n232_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n225_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n218_), .A2(new_n236_), .A3(new_n235_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n230_), .B1(new_n240_), .B2(new_n229_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n213_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n229_), .B1(new_n237_), .B2(new_n232_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n230_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n245_), .A2(new_n212_), .A3(new_n225_), .A4(new_n238_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(KEYINPUT12), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n225_), .A3(new_n238_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT12), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(new_n213_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n204_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n242_), .A2(new_n246_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n204_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G120gat), .B(G148gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G176gat), .B(G204gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n255_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n252_), .A2(new_n254_), .A3(new_n260_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT13), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n263_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT13), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT67), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT72), .ZN(new_n273_));
  XOR2_X1   g072(.A(G127gat), .B(G155gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G183gat), .B(G211gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT17), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G231gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n212_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G8gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT14), .ZN(new_n283_));
  OR2_X1    g082(.A1(KEYINPUT70), .A2(G1gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(KEYINPUT70), .A2(G1gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n283_), .B1(new_n286_), .B2(G8gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(G15gat), .B(G22gat), .Z(new_n288_));
  OAI21_X1  g087(.A(new_n282_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  INV_X1    g089(.A(G8gat), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n290_), .B(new_n281_), .C1(new_n292_), .C2(new_n283_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n280_), .B(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n278_), .A2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n277_), .A2(KEYINPUT17), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n278_), .A3(new_n296_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n297_), .A2(new_n299_), .A3(KEYINPUT73), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT73), .B1(new_n299_), .B2(new_n297_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT69), .B(KEYINPUT37), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G29gat), .B(G36gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(G43gat), .B(G50gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT15), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n248_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G232gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT34), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n315_), .A2(KEYINPUT35), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n311_), .B1(new_n308_), .B2(new_n248_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G190gat), .B(G218gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G134gat), .B(G162gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n317_), .A2(new_n318_), .B1(KEYINPUT36), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n318_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n315_), .A2(KEYINPUT35), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n315_), .A2(KEYINPUT35), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n323_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n321_), .A2(KEYINPUT36), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n322_), .B2(new_n327_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n305_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n322_), .A2(new_n327_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n328_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n330_), .A3(new_n304_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n271_), .A2(new_n303_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n308_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n294_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G229gat), .A2(G233gat), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n310_), .A2(new_n295_), .A3(KEYINPUT76), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT76), .B1(new_n310_), .B2(new_n295_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n340_), .B(new_n341_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n289_), .A2(new_n308_), .A3(new_n293_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n308_), .B1(new_n293_), .B2(new_n289_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n289_), .A2(new_n308_), .A3(new_n293_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n340_), .A2(KEYINPUT74), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n341_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT75), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354_));
  AOI211_X1 g153(.A(new_n354_), .B(new_n341_), .C1(new_n348_), .C2(new_n350_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n344_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G113gat), .B(G141gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT77), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G169gat), .B(G197gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n360_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n344_), .B(new_n362_), .C1(new_n353_), .C2(new_n355_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT78), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G211gat), .B(G218gat), .Z(new_n370_));
  OR2_X1    g169(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n371_));
  INV_X1    g170(.A(G204gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT21), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(G197gat), .B2(G204gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n370_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n371_), .A2(G204gat), .A3(new_n373_), .ZN(new_n378_));
  INV_X1    g177(.A(G197gat), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n379_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT90), .B1(new_n379_), .B2(G204gat), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n378_), .A2(new_n380_), .A3(new_n375_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n370_), .A2(KEYINPUT21), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n378_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G141gat), .A2(G148gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(KEYINPUT1), .B2(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n392_), .A2(KEYINPUT1), .ZN(new_n394_));
  AOI211_X1 g193(.A(new_n388_), .B(new_n390_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT2), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n389_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT85), .B(KEYINPUT3), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT86), .B1(new_n402_), .B2(new_n388_), .ZN(new_n403_));
  AND2_X1   g202(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n404_));
  NOR2_X1   g203(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n405_));
  OAI211_X1 g204(.A(KEYINPUT86), .B(new_n388_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n401_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n392_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(new_n391_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n395_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n387_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT88), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n414_), .A2(KEYINPUT88), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n387_), .A2(KEYINPUT91), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n382_), .A2(new_n377_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n393_), .A2(new_n394_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n390_), .A2(new_n388_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n388_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n400_), .B1(new_n425_), .B2(new_n406_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n410_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n422_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n419_), .B1(new_n428_), .B2(KEYINPUT29), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n416_), .A2(new_n415_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT91), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n430_), .B1(new_n419_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G78gat), .B(G106gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n418_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n418_), .B2(new_n433_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n440_));
  OR3_X1    g239(.A1(new_n428_), .A2(KEYINPUT29), .A3(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G22gat), .B(G50gat), .Z(new_n442_));
  OAI21_X1  g241(.A(new_n440_), .B1(new_n428_), .B2(KEYINPUT29), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n442_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT92), .B1(new_n439_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT93), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n438_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n438_), .A2(new_n448_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n449_), .A2(new_n446_), .A3(new_n436_), .A4(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n444_), .A2(new_n445_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT92), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n452_), .B(new_n453_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n447_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G169gat), .ZN(new_n456_));
  INV_X1    g255(.A(G176gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(KEYINPUT24), .A3(new_n459_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n458_), .A2(KEYINPUT24), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G183gat), .A2(G190gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT81), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(G183gat), .A3(G190gat), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT23), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT23), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(G183gat), .B2(G190gat), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n460_), .B(new_n461_), .C1(new_n466_), .C2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(G190gat), .ZN(new_n471_));
  INV_X1    g270(.A(G190gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(KEYINPUT80), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT26), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT25), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT25), .ZN(new_n480_));
  INV_X1    g279(.A(G183gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n474_), .A2(new_n476_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n469_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n456_), .A2(KEYINPUT22), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT22), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G169gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n487_), .A3(new_n457_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT82), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT22), .B(G169gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT82), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n457_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n489_), .A2(new_n492_), .A3(new_n459_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT83), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n462_), .A2(new_n467_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n463_), .A2(new_n465_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(KEYINPUT23), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n477_), .A2(new_n478_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT80), .B(G190gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n493_), .A2(new_n494_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n459_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n503_), .B1(new_n488_), .B2(KEYINPUT82), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT83), .A3(new_n492_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n484_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT97), .B1(new_n506_), .B2(new_n419_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n493_), .A2(new_n494_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n498_), .A2(new_n501_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n484_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT97), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n387_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n507_), .A2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(new_n475_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n519_), .A2(new_n520_), .A3(KEYINPUT94), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT94), .ZN(new_n522_));
  NAND2_X1  g321(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n482_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n518_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n460_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT94), .B1(new_n519_), .B2(new_n520_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n482_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n517_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n460_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT95), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n498_), .A2(new_n461_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n527_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT96), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n468_), .B1(new_n497_), .B2(new_n467_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G183gat), .A2(G190gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OAI221_X1 g337(.A(KEYINPUT96), .B1(G183gat), .B2(G190gat), .C1(new_n466_), .C2(new_n468_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n503_), .B1(new_n490_), .B2(new_n457_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n534_), .A2(new_n419_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G226gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT19), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n542_), .A2(KEYINPUT20), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n515_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n534_), .A2(new_n541_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n387_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n510_), .A2(new_n511_), .A3(new_n419_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(KEYINPUT20), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n544_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G8gat), .B(G36gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT18), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G64gat), .B(G92gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT32), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n547_), .A2(new_n552_), .A3(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G1gat), .B(G29gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(G85gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT0), .B(G57gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  XNOR2_X1  g361(.A(G127gat), .B(G134gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G113gat), .B(G120gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n411_), .B2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n422_), .B(new_n567_), .C1(new_n426_), .C2(new_n427_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(new_n565_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT4), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G225gat), .A2(G233gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n565_), .A2(KEYINPUT4), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n428_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT100), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT100), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n428_), .A2(new_n577_), .A3(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n571_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n572_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n562_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n428_), .A2(new_n577_), .A3(new_n574_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n577_), .B1(new_n428_), .B2(new_n574_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n573_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT4), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n411_), .A2(new_n567_), .A3(new_n566_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n569_), .A2(new_n565_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n586_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n581_), .B(new_n562_), .C1(new_n585_), .C2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n558_), .B1(new_n582_), .B2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n542_), .A2(KEYINPUT20), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n513_), .B1(new_n512_), .B2(new_n387_), .ZN(new_n594_));
  AOI211_X1 g393(.A(KEYINPUT97), .B(new_n419_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n593_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n544_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n551_), .A2(new_n544_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n557_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT102), .B1(new_n592_), .B2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n545_), .B1(new_n515_), .B2(new_n593_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n551_), .A2(new_n544_), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT32), .B(new_n556_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT102), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n581_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n562_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n590_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n603_), .A2(new_n604_), .A3(new_n608_), .A4(new_n558_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n600_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n547_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT98), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n547_), .A2(new_n552_), .A3(new_n613_), .A4(new_n556_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n547_), .A2(new_n552_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n556_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n591_), .A2(KEYINPUT33), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n571_), .A2(new_n572_), .A3(new_n579_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n568_), .A2(new_n570_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n621_), .A2(KEYINPUT101), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n573_), .B1(new_n621_), .B2(KEYINPUT101), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n620_), .B(new_n606_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n590_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n619_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n618_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n455_), .B1(new_n610_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT27), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n616_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n611_), .A2(KEYINPUT27), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n618_), .A2(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n608_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n447_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n629_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G71gat), .B(G99gat), .ZN(new_n638_));
  INV_X1    g437(.A(G43gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT30), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G227gat), .A2(G233gat), .ZN(new_n642_));
  INV_X1    g441(.A(G15gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n641_), .B(new_n644_), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n506_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT31), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(new_n506_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n646_), .A2(KEYINPUT84), .A3(new_n647_), .A4(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(KEYINPUT84), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT31), .B1(new_n651_), .B2(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n565_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n650_), .A2(new_n566_), .A3(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n637_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n654_), .A2(new_n634_), .A3(new_n655_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n633_), .A2(KEYINPUT103), .A3(new_n455_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT103), .B1(new_n633_), .B2(new_n455_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n369_), .B1(new_n657_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n338_), .A2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n608_), .B(KEYINPUT104), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT105), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT38), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n331_), .A2(new_n332_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n657_), .B2(new_n662_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n299_), .A2(new_n297_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n269_), .A2(new_n365_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G1gat), .B1(new_n675_), .B2(new_n634_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n668_), .A2(KEYINPUT38), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n669_), .A2(new_n676_), .A3(new_n677_), .ZN(G1324gat));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n679_));
  NOR4_X1   g478(.A1(new_n269_), .A2(new_n633_), .A3(new_n365_), .A4(new_n672_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n670_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n618_), .A2(new_n630_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n632_), .A2(new_n631_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n455_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n633_), .A2(KEYINPUT103), .A3(new_n455_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n658_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n654_), .A2(new_n655_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n629_), .B2(new_n636_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n680_), .B(new_n681_), .C1(new_n688_), .C2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(KEYINPUT106), .A3(G8gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT106), .B1(new_n691_), .B2(G8gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n679_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n694_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(KEYINPUT107), .A3(new_n692_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n697_), .A3(KEYINPUT39), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT39), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n679_), .B(new_n699_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n664_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n633_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n291_), .A3(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n698_), .A2(new_n700_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT40), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n698_), .A2(KEYINPUT40), .A3(new_n700_), .A4(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1325gat));
  OAI21_X1  g507(.A(G15gat), .B1(new_n675_), .B2(new_n656_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT41), .Z(new_n710_));
  NAND3_X1  g509(.A1(new_n701_), .A2(new_n643_), .A3(new_n689_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1326gat));
  OAI21_X1  g511(.A(G22gat), .B1(new_n675_), .B2(new_n455_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT42), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n455_), .A2(G22gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n664_), .B2(new_n715_), .ZN(G1327gat));
  NAND2_X1  g515(.A1(new_n303_), .A2(new_n670_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n269_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n663_), .A2(new_n718_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n719_), .A2(G29gat), .A3(new_n634_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n333_), .A2(new_n336_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT109), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n723_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n657_), .A2(new_n662_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n722_), .A2(KEYINPUT43), .ZN(new_n727_));
  AOI22_X1  g526(.A1(new_n724_), .A2(new_n725_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n674_), .A2(new_n303_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n721_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n729_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n725_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n726_), .B2(new_n723_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n727_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n657_), .B2(new_n662_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT44), .B(new_n731_), .C1(new_n733_), .C2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n730_), .A2(new_n665_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n720_), .B1(new_n737_), .B2(G29gat), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT110), .B(new_n720_), .C1(new_n737_), .C2(G29gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1328gat));
  NAND3_X1  g541(.A1(new_n730_), .A2(new_n702_), .A3(new_n736_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G36gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n633_), .A2(G36gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n663_), .A2(new_n718_), .A3(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT45), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n744_), .A2(KEYINPUT46), .A3(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1329gat));
  NAND4_X1  g551(.A1(new_n730_), .A2(G43gat), .A3(new_n736_), .A4(new_n689_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n639_), .B1(new_n719_), .B2(new_n656_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g555(.A1(new_n730_), .A2(new_n635_), .A3(new_n736_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(G50gat), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n455_), .A2(G50gat), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT111), .Z(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n719_), .B2(new_n760_), .ZN(G1331gat));
  AOI21_X1  g560(.A(new_n364_), .B1(new_n657_), .B2(new_n662_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n762_), .A2(new_n269_), .A3(new_n302_), .A4(new_n722_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G57gat), .B1(new_n764_), .B2(new_n665_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n302_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n270_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n671_), .A2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(KEYINPUT112), .B(G57gat), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n768_), .A2(new_n634_), .A3(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n765_), .A2(new_n770_), .ZN(G1332gat));
  OAI21_X1  g570(.A(G64gat), .B1(new_n768_), .B2(new_n633_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT48), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n633_), .A2(G64gat), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT113), .Z(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n763_), .B2(new_n775_), .ZN(G1333gat));
  OR3_X1    g575(.A1(new_n763_), .A2(G71gat), .A3(new_n656_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n671_), .A2(new_n689_), .A3(new_n767_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(G71gat), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n778_), .B2(G71gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n777_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT114), .ZN(G1334gat));
  OAI21_X1  g583(.A(G78gat), .B1(new_n768_), .B2(new_n455_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT50), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n455_), .A2(G78gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n763_), .B2(new_n787_), .ZN(G1335gat));
  AND3_X1   g587(.A1(new_n303_), .A2(new_n365_), .A3(new_n269_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n634_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n762_), .A2(new_n271_), .A3(new_n303_), .A4(new_n670_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n221_), .A3(new_n665_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(G1336gat));
  OAI21_X1  g594(.A(G92gat), .B1(new_n790_), .B2(new_n633_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n222_), .A3(new_n702_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1337gat));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n800_));
  OAI21_X1  g599(.A(G99gat), .B1(new_n790_), .B2(new_n656_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n793_), .A2(new_n689_), .A3(new_n214_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(G1338gat));
  NAND3_X1  g604(.A1(new_n793_), .A2(new_n215_), .A3(new_n635_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n635_), .B(new_n789_), .C1(new_n733_), .C2(new_n735_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n215_), .B1(KEYINPUT116), .B2(KEYINPUT52), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n806_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT53), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n814_), .B(new_n806_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(G1339gat));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n340_), .B(new_n352_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n351_), .A2(new_n341_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n360_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n363_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n363_), .A2(KEYINPUT120), .A3(new_n820_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n264_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT119), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n247_), .A2(new_n204_), .A3(new_n250_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n829_), .A2(new_n251_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n251_), .A2(new_n830_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n261_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n827_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n252_), .A2(KEYINPUT55), .A3(new_n828_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n260_), .B1(new_n251_), .B2(new_n830_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n835_), .A2(KEYINPUT119), .A3(new_n826_), .A4(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n263_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n838_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n364_), .A2(new_n263_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT118), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n825_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n817_), .B1(new_n845_), .B2(new_n670_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n823_), .A2(new_n824_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n266_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n364_), .A2(new_n841_), .A3(new_n263_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n834_), .A2(new_n837_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n840_), .A2(new_n841_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n848_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(KEYINPUT57), .A3(new_n681_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n831_), .A2(new_n833_), .A3(KEYINPUT56), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n826_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n855_), .A2(new_n839_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n847_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n857_), .A2(new_n847_), .A3(KEYINPUT58), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n337_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n846_), .A2(new_n854_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n672_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n333_), .A2(new_n265_), .A3(new_n336_), .A4(new_n268_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n866_), .A2(new_n369_), .A3(new_n302_), .A4(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n867_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n766_), .B2(new_n865_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n864_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n660_), .A2(new_n661_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n689_), .A2(new_n665_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(G113gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n878_), .A3(new_n364_), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT121), .B1(new_n863_), .B2(new_n303_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n863_), .A2(KEYINPUT121), .A3(new_n303_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n871_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n875_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(KEYINPUT59), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n871_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n672_), .B2(new_n863_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT59), .B1(new_n889_), .B2(new_n884_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n887_), .A2(new_n891_), .A3(new_n369_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n879_), .B1(new_n892_), .B2(new_n878_), .ZN(G1340gat));
  AND3_X1   g692(.A1(new_n863_), .A2(KEYINPUT121), .A3(new_n303_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n894_), .A2(new_n880_), .A3(new_n888_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n885_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n890_), .B(new_n271_), .C1(new_n895_), .C2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT123), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n886_), .A2(new_n899_), .A3(new_n271_), .A4(new_n890_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n898_), .A2(G120gat), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n902_));
  AOI21_X1  g701(.A(KEYINPUT122), .B1(new_n902_), .B2(G120gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(G120gat), .B1(new_n269_), .B2(new_n902_), .ZN(new_n904_));
  MUX2_X1   g703(.A(new_n903_), .B(KEYINPUT122), .S(new_n904_), .Z(new_n905_));
  NAND2_X1  g704(.A1(new_n877_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n901_), .A2(new_n906_), .ZN(G1341gat));
  NOR2_X1   g706(.A1(new_n876_), .A2(new_n303_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n908_), .A2(new_n909_), .A3(G127gat), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n886_), .A2(G127gat), .A3(new_n673_), .A4(new_n890_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n908_), .B2(G127gat), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(G1342gat));
  INV_X1    g712(.A(G134gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n877_), .A2(new_n914_), .A3(new_n670_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n887_), .A2(new_n891_), .A3(new_n722_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n914_), .ZN(G1343gat));
  NAND4_X1  g716(.A1(new_n656_), .A2(new_n635_), .A3(new_n633_), .A4(new_n665_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT125), .Z(new_n919_));
  NAND2_X1  g718(.A1(new_n872_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n365_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT126), .B(G141gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1344gat));
  INV_X1    g722(.A(new_n920_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n271_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g725(.A1(new_n920_), .A2(new_n303_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT61), .B(G155gat), .Z(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1346gat));
  AOI21_X1  g728(.A(G162gat), .B1(new_n924_), .B2(new_n670_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n723_), .A2(G162gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n924_), .B2(new_n931_), .ZN(G1347gat));
  OR3_X1    g731(.A1(new_n656_), .A2(new_n633_), .A3(new_n665_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n635_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n883_), .A2(new_n934_), .ZN(new_n935_));
  OAI21_X1  g734(.A(G169gat), .B1(new_n935_), .B2(new_n365_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n935_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n939_), .A2(new_n490_), .A3(new_n364_), .ZN(new_n940_));
  OAI211_X1 g739(.A(KEYINPUT62), .B(G169gat), .C1(new_n935_), .C2(new_n365_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n938_), .A2(new_n940_), .A3(new_n941_), .ZN(G1348gat));
  AOI21_X1  g741(.A(G176gat), .B1(new_n939_), .B2(new_n269_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n889_), .A2(new_n635_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n933_), .A2(new_n270_), .A3(new_n457_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n943_), .B1(new_n944_), .B2(new_n945_), .ZN(G1349gat));
  NOR3_X1   g745(.A1(new_n672_), .A2(new_n524_), .A3(new_n521_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n933_), .A2(new_n303_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n944_), .A2(new_n948_), .ZN(new_n949_));
  AOI22_X1  g748(.A1(new_n939_), .A2(new_n947_), .B1(new_n499_), .B2(new_n949_), .ZN(G1350gat));
  OAI21_X1  g749(.A(G190gat), .B1(new_n935_), .B2(new_n722_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n670_), .A2(new_n518_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n935_), .B2(new_n952_), .ZN(G1351gat));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n656_), .A2(new_n634_), .A3(new_n702_), .A4(new_n635_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n889_), .B2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n955_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n872_), .A2(KEYINPUT127), .A3(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n956_), .A2(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(new_n364_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g760(.A1(new_n959_), .A2(new_n271_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g762(.A(KEYINPUT63), .B(G211gat), .C1(new_n959_), .C2(new_n673_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(KEYINPUT63), .B(G211gat), .ZN(new_n965_));
  AOI211_X1 g764(.A(new_n672_), .B(new_n965_), .C1(new_n956_), .C2(new_n958_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n964_), .A2(new_n966_), .ZN(G1354gat));
  INV_X1    g766(.A(G218gat), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n959_), .A2(new_n968_), .A3(new_n670_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n722_), .B1(new_n956_), .B2(new_n958_), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n969_), .B1(new_n968_), .B2(new_n970_), .ZN(G1355gat));
endmodule


