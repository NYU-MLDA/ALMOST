//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n950_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n214_), .A2(new_n217_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G85gat), .B(G92gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(KEYINPUT8), .A3(new_n221_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT10), .B(G99gat), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n213_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(KEYINPUT9), .ZN(new_n229_));
  INV_X1    g028(.A(G85gat), .ZN(new_n230_));
  INV_X1    g029(.A(G92gat), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT9), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n217_), .A2(new_n218_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n210_), .B1(new_n226_), .B2(new_n234_), .ZN(new_n235_));
  AND4_X1   g034(.A1(new_n210_), .A2(new_n234_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n236_));
  OAI211_X1 g035(.A(KEYINPUT12), .B(new_n209_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n208_), .A2(new_n225_), .A3(new_n234_), .A4(new_n224_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n239_), .A2(KEYINPUT12), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(KEYINPUT12), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n226_), .A2(new_n234_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n209_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G230gat), .A2(G233gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n237_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n238_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(G230gat), .A3(G233gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G120gat), .B(G148gat), .ZN(new_n251_));
  INV_X1    g050(.A(G204gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT5), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G176gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n250_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT13), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(KEYINPUT67), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n256_), .B(KEYINPUT66), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT67), .B(KEYINPUT13), .Z(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G15gat), .B(G22gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT69), .B(G8gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT14), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G1gat), .ZN(new_n270_));
  INV_X1    g069(.A(G1gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n266_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G8gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G29gat), .B(G36gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(G43gat), .ZN(new_n277_));
  INV_X1    g076(.A(G50gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT72), .ZN(new_n281_));
  INV_X1    g080(.A(new_n275_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n277_), .B(G50gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n281_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G229gat), .A2(G233gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n280_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n279_), .A2(KEYINPUT15), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT15), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n283_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n282_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n286_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n288_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G113gat), .B(G141gat), .ZN(new_n297_));
  INV_X1    g096(.A(G169gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G197gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n288_), .A2(new_n295_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n265_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G176gat), .ZN(new_n308_));
  AND2_X1   g107(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317_));
  NAND3_X1  g116(.A1(KEYINPUT75), .A2(G183gat), .A3(G190gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(KEYINPUT74), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT23), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n322_), .A3(new_n314_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n313_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n317_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n314_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(KEYINPUT89), .A2(KEYINPUT24), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n298_), .A2(new_n308_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(KEYINPUT89), .A2(KEYINPUT24), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n312_), .A4(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n333_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n335_), .B1(new_n336_), .B2(new_n330_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n329_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G190gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT25), .B(G183gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n326_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n252_), .A2(G197gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n300_), .A2(G204gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT83), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(G197gat), .B2(new_n252_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT21), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n346_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .A4(KEYINPUT21), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G211gat), .A2(G218gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G211gat), .A2(G218gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n352_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(G211gat), .A2(G218gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(KEYINPUT84), .A3(new_n353_), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n350_), .A2(new_n351_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT86), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n349_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n361_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n359_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n356_), .A2(new_n358_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n351_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT83), .B1(new_n300_), .B2(G204gat), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n366_), .A2(KEYINPUT21), .B1(new_n344_), .B2(new_n345_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n364_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n361_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT86), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n343_), .B1(new_n363_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n325_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n313_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT73), .ZN(new_n375_));
  INV_X1    g174(.A(G183gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(KEYINPUT25), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n377_), .B(new_n340_), .C1(new_n341_), .C2(new_n375_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n379_));
  AND2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(new_n335_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n381_), .B2(KEYINPUT24), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(new_n324_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n374_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n368_), .A2(new_n369_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n384_), .A2(KEYINPUT91), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT91), .B1(new_n384_), .B2(new_n385_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n371_), .B(KEYINPUT20), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT19), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n388_), .A2(KEYINPUT95), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT95), .B1(new_n388_), .B2(new_n390_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n393_));
  INV_X1    g192(.A(new_n384_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n385_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT90), .B1(new_n343_), .B2(new_n395_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT90), .ZN(new_n398_));
  INV_X1    g197(.A(new_n342_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n329_), .A2(new_n399_), .A3(new_n338_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n398_), .B(new_n385_), .C1(new_n400_), .C2(new_n326_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n396_), .A2(new_n397_), .A3(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n390_), .B(KEYINPUT88), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n391_), .A2(new_n392_), .A3(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT96), .B1(new_n406_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n402_), .A2(new_n404_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n393_), .B1(new_n343_), .B2(new_n395_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n390_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n414_), .B(new_n415_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n413_), .A2(new_n416_), .A3(new_n411_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n388_), .A2(new_n390_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT95), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n405_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n388_), .A2(KEYINPUT95), .A3(new_n390_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT96), .ZN(new_n425_));
  INV_X1    g224(.A(new_n411_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n412_), .A2(KEYINPUT27), .A3(new_n418_), .A4(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT30), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n374_), .A2(new_n430_), .A3(new_n383_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n374_), .B2(new_n383_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n383_), .ZN(new_n434_));
  AND3_X1   g233(.A1(KEYINPUT75), .A2(G183gat), .A3(G190gat), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT75), .B1(G183gat), .B2(G190gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT23), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT74), .B(KEYINPUT23), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n314_), .B2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n313_), .B1(new_n439_), .B2(new_n325_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT30), .B1(new_n434_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n429_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n374_), .A2(new_n430_), .A3(new_n383_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445_));
  INV_X1    g244(.A(G15gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(G43gat), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n433_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n448_), .B1(new_n433_), .B2(new_n444_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT77), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n448_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n431_), .A2(new_n432_), .A3(new_n429_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n442_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT77), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n433_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(G127gat), .A2(G134gat), .ZN(new_n459_));
  INV_X1    g258(.A(G113gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G127gat), .A2(G134gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(G127gat), .A2(G134gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G127gat), .A2(G134gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(G113gat), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n462_), .A2(new_n465_), .A3(G120gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(G120gat), .B1(new_n462_), .B2(new_n465_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n451_), .A2(new_n458_), .A3(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(KEYINPUT77), .B(new_n470_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G228gat), .A2(G233gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n475_), .B(KEYINPUT81), .Z(new_n476_));
  OAI21_X1  g275(.A(new_n360_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n368_), .A2(KEYINPUT86), .A3(new_n369_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT2), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT78), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n482_), .A3(new_n480_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT3), .ZN(new_n487_));
  INV_X1    g286(.A(G141gat), .ZN(new_n488_));
  INV_X1    g287(.A(G148gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .A4(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(G155gat), .A2(G162gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G155gat), .A2(G162gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT1), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n494_), .A2(new_n495_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n492_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n491_), .A2(new_n494_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT85), .B(KEYINPUT29), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n476_), .B1(new_n479_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT29), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT80), .B1(new_n498_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n488_), .A2(new_n489_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G155gat), .B(G162gat), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n497_), .B(new_n504_), .C1(KEYINPUT1), .C2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n490_), .A2(new_n486_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n481_), .A2(new_n482_), .A3(new_n480_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n483_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n506_), .B1(new_n509_), .B2(new_n505_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT80), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT29), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n476_), .B(KEYINPUT82), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n503_), .A2(new_n385_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n501_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G78gat), .B(G106gat), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n501_), .A2(new_n516_), .A3(new_n514_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n501_), .A2(new_n514_), .A3(new_n520_), .A4(new_n516_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT79), .B(KEYINPUT28), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n510_), .B2(KEYINPUT29), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n498_), .A2(new_n502_), .A3(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G22gat), .B(G50gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n518_), .A2(new_n519_), .B1(new_n521_), .B2(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n501_), .A2(new_n516_), .A3(new_n514_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n516_), .B1(new_n501_), .B2(new_n514_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n523_), .A2(new_n525_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n526_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(KEYINPUT87), .A3(new_n527_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n532_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n531_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n474_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n518_), .A2(KEYINPUT87), .A3(new_n519_), .A4(new_n530_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n532_), .A2(new_n533_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n521_), .A2(new_n530_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(new_n473_), .A3(new_n472_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT27), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n411_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n417_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT97), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT97), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n551_), .B(new_n547_), .C1(new_n417_), .C2(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n498_), .A2(new_n468_), .A3(KEYINPUT93), .ZN(new_n554_));
  OAI211_X1 g353(.A(KEYINPUT93), .B(new_n506_), .C1(new_n509_), .C2(new_n505_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n467_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n462_), .A2(new_n465_), .A3(G120gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G225gat), .A2(G233gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n498_), .A2(new_n468_), .A3(KEYINPUT4), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n559_), .A3(KEYINPUT4), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT94), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n554_), .A2(new_n559_), .A3(new_n566_), .A4(KEYINPUT4), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n563_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n562_), .B1(new_n568_), .B2(new_n561_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT0), .B(G57gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G85gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(G1gat), .B(G29gat), .Z(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n573_), .B(new_n562_), .C1(new_n568_), .C2(new_n561_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n428_), .A2(new_n546_), .A3(new_n553_), .A4(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n568_), .A2(new_n561_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n582_), .B(new_n573_), .C1(new_n561_), .C2(new_n560_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n417_), .A2(new_n548_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n569_), .A2(KEYINPUT33), .A3(new_n574_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n581_), .A2(new_n583_), .A3(new_n584_), .A4(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n411_), .A2(KEYINPUT32), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n424_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n411_), .A2(KEYINPUT32), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n413_), .A2(new_n416_), .A3(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n577_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n474_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n539_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n579_), .A2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n307_), .A2(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n235_), .A2(new_n236_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n293_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT34), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT35), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n279_), .A2(new_n234_), .A3(new_n226_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n599_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n602_), .A2(new_n603_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n599_), .A2(KEYINPUT35), .A3(new_n601_), .A4(new_n605_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(G134gat), .ZN(new_n613_));
  INV_X1    g412(.A(G162gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  AOI22_X1  g414(.A1(new_n609_), .A2(new_n610_), .B1(new_n611_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n615_), .B(KEYINPUT36), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n609_), .A2(new_n619_), .A3(new_n610_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT37), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n617_), .A2(new_n620_), .A3(KEYINPUT68), .A4(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(KEYINPUT68), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(KEYINPUT68), .ZN(new_n624_));
  INV_X1    g423(.A(new_n620_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n623_), .B(new_n624_), .C1(new_n625_), .C2(new_n616_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n275_), .B(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n208_), .B(KEYINPUT70), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(G127gat), .B(G155gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT71), .B(KEYINPUT16), .Z(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT17), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n631_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n636_), .A2(KEYINPUT17), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n639_), .B1(new_n642_), .B2(new_n631_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n627_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n597_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n271_), .A3(new_n577_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT38), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n625_), .A2(new_n616_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI211_X1 g449(.A(new_n643_), .B(new_n650_), .C1(new_n579_), .C2(new_n595_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n307_), .A2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT98), .Z(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n578_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n648_), .A2(new_n654_), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n428_), .A2(new_n553_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G8gat), .B1(new_n652_), .B2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT39), .Z(new_n659_));
  NOR3_X1   g458(.A1(new_n645_), .A2(new_n267_), .A3(new_n657_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g461(.A(G15gat), .B1(new_n653_), .B2(new_n474_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT41), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n646_), .A2(new_n446_), .A3(new_n593_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1326gat));
  XNOR2_X1  g465(.A(new_n544_), .B(KEYINPUT99), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G22gat), .B1(new_n653_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT42), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(G22gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT100), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n645_), .B2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n596_), .A2(new_n674_), .A3(new_n627_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n627_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n596_), .B2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n579_), .A2(new_n595_), .A3(KEYINPUT101), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT102), .B(new_n674_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n596_), .A2(new_n677_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n627_), .A3(new_n679_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n683_), .B2(KEYINPUT43), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n675_), .B1(new_n680_), .B2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n307_), .A3(new_n643_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n687_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n685_), .A2(new_n307_), .A3(new_n643_), .A4(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n578_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n643_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n649_), .A2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n597_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(G29gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n577_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n692_), .A2(new_n697_), .ZN(G1328gat));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(new_n699_), .A3(new_n656_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT45), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n691_), .A2(new_n657_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(new_n699_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(KEYINPUT46), .B(new_n701_), .C1(new_n702_), .C2(new_n699_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  AOI21_X1  g506(.A(G43gat), .B1(new_n695_), .B2(new_n593_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT104), .Z(new_n709_));
  NAND4_X1  g508(.A1(new_n688_), .A2(G43gat), .A3(new_n593_), .A4(new_n690_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT47), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n713_), .A3(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1330gat));
  OAI21_X1  g514(.A(G50gat), .B1(new_n691_), .B2(new_n544_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n695_), .A2(new_n278_), .A3(new_n667_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n264_), .A2(new_n305_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(new_n651_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n578_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n596_), .A2(new_n306_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT105), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(new_n264_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n644_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n727_), .A2(KEYINPUT106), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(KEYINPUT106), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n577_), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n723_), .B1(new_n730_), .B2(new_n722_), .ZN(G1332gat));
  INV_X1    g530(.A(G64gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n720_), .B2(new_n656_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT48), .Z(new_n734_));
  NAND2_X1  g533(.A1(new_n656_), .A2(new_n732_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n727_), .B2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n721_), .B2(new_n474_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT107), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT49), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n474_), .A2(G71gat), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n740_), .A2(new_n741_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n726_), .A2(new_n644_), .A3(new_n742_), .A4(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n739_), .A2(new_n744_), .ZN(G1334gat));
  INV_X1    g544(.A(G78gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n720_), .B2(new_n667_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT50), .Z(new_n748_));
  NAND2_X1  g547(.A1(new_n667_), .A2(new_n746_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n727_), .B2(new_n749_), .ZN(G1335gat));
  AND2_X1   g549(.A1(new_n685_), .A2(KEYINPUT109), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n685_), .A2(KEYINPUT109), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n719_), .A2(new_n643_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(G85gat), .A3(new_n577_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n726_), .A2(new_n694_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n230_), .B1(new_n756_), .B2(new_n578_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1336gat));
  NAND3_X1  g557(.A1(new_n754_), .A2(G92gat), .A3(new_n656_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n231_), .B1(new_n756_), .B2(new_n657_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1337gat));
  NAND2_X1  g560(.A1(new_n754_), .A2(new_n593_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G99gat), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n726_), .A2(new_n227_), .A3(new_n593_), .A4(new_n694_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT51), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(new_n767_), .A3(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1338gat));
  INV_X1    g568(.A(new_n675_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n579_), .A2(new_n595_), .A3(KEYINPUT101), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT101), .B1(new_n579_), .B2(new_n595_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n676_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT102), .B1(new_n773_), .B2(new_n674_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n683_), .A2(new_n681_), .A3(KEYINPUT43), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n770_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n753_), .A2(new_n544_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT110), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n685_), .A2(new_n780_), .A3(new_n777_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(G106gat), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT111), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n779_), .A2(new_n781_), .A3(new_n784_), .A4(G106gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(KEYINPUT52), .A3(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n726_), .A2(new_n213_), .A3(new_n539_), .A4(new_n694_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n782_), .A2(KEYINPUT111), .A3(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT53), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n786_), .A2(new_n792_), .A3(new_n787_), .A4(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1339gat));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n285_), .A2(new_n286_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n294_), .A2(new_n287_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n301_), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n304_), .A3(KEYINPUT116), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n304_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n258_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n246_), .B1(new_n237_), .B2(new_n245_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n247_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n237_), .A2(new_n245_), .A3(KEYINPUT55), .A4(new_n246_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n255_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n808_), .A2(KEYINPUT114), .A3(new_n255_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n810_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n811_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n813_), .A2(KEYINPUT115), .A3(new_n810_), .A4(new_n814_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n306_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n250_), .A2(new_n255_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n803_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n795_), .B1(new_n822_), .B2(new_n650_), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n306_), .B(new_n820_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT57), .B(new_n649_), .C1(new_n824_), .C2(new_n803_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n802_), .A2(new_n799_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n809_), .B(new_n810_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n821_), .A3(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT58), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n627_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n823_), .A2(new_n825_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n643_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n305_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n644_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n835_), .B2(new_n644_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n834_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(new_n644_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT112), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n837_), .A3(new_n833_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n840_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n832_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n656_), .A2(new_n578_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n845_), .A2(new_n593_), .A3(new_n544_), .A4(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G113gat), .B1(new_n848_), .B2(new_n305_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(KEYINPUT118), .A2(G113gat), .ZN(new_n850_));
  AND2_X1   g649(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n847_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n850_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G113gat), .B1(new_n306_), .B2(KEYINPUT118), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n849_), .B1(new_n856_), .B2(new_n857_), .ZN(G1340gat));
  AOI21_X1  g657(.A(new_n264_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n859_));
  INV_X1    g658(.A(G120gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(KEYINPUT60), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n847_), .A2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n264_), .B2(KEYINPUT60), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT119), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865_));
  INV_X1    g664(.A(new_n863_), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n847_), .A2(new_n865_), .A3(new_n866_), .A4(new_n861_), .ZN(new_n867_));
  OAI22_X1  g666(.A1(new_n859_), .A2(new_n860_), .B1(new_n864_), .B2(new_n867_), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n848_), .B2(new_n693_), .ZN(new_n869_));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n871_), .B2(new_n693_), .ZN(G1342gat));
  AOI21_X1  g671(.A(G134gat), .B1(new_n848_), .B2(new_n650_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n676_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(G134gat), .ZN(G1343gat));
  XNOR2_X1  g674(.A(KEYINPUT121), .B(G141gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n540_), .B1(new_n832_), .B2(new_n844_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n846_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n877_), .A2(KEYINPUT120), .A3(new_n846_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n876_), .B1(new_n882_), .B2(new_n305_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n840_), .A2(new_n843_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n643_), .B2(new_n831_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n846_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n885_), .A2(new_n879_), .A3(new_n540_), .A4(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT120), .B1(new_n877_), .B2(new_n846_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n305_), .B(new_n876_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n883_), .A2(new_n890_), .ZN(G1344gat));
  XNOR2_X1  g690(.A(KEYINPUT122), .B(G148gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n882_), .B2(new_n265_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n265_), .B(new_n892_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1345gat));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n882_), .B2(new_n693_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n693_), .B(new_n897_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1346gat));
  NAND2_X1  g700(.A1(new_n882_), .A2(new_n650_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n627_), .A2(G162gat), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT123), .Z(new_n904_));
  AOI22_X1  g703(.A1(new_n902_), .A2(new_n614_), .B1(new_n882_), .B2(new_n904_), .ZN(G1347gat));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n657_), .A2(new_n577_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n474_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n845_), .A2(new_n305_), .A3(new_n668_), .A4(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n911_), .A3(G169gat), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n910_), .B2(G169gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n906_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n909_), .ZN(new_n916_));
  NOR4_X1   g715(.A1(new_n885_), .A2(new_n306_), .A3(new_n667_), .A4(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT124), .B1(new_n917_), .B2(new_n298_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(KEYINPUT62), .A3(new_n912_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n917_), .B1(new_n310_), .B2(new_n309_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n915_), .A2(new_n919_), .A3(new_n920_), .ZN(G1348gat));
  NOR3_X1   g720(.A1(new_n885_), .A2(new_n667_), .A3(new_n916_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n922_), .A2(new_n308_), .A3(new_n265_), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n885_), .A2(new_n264_), .A3(new_n539_), .A4(new_n916_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n308_), .B2(new_n924_), .ZN(G1349gat));
  INV_X1    g724(.A(new_n922_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n926_), .A2(new_n643_), .A3(new_n341_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n845_), .A2(new_n693_), .A3(new_n544_), .A4(new_n909_), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT125), .Z(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n929_), .B2(new_n376_), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n926_), .B2(new_n676_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n922_), .A2(new_n340_), .A3(new_n650_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1351gat));
  NAND2_X1  g732(.A1(new_n877_), .A2(new_n907_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n306_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n300_), .ZN(G1352gat));
  NOR2_X1   g735(.A1(new_n934_), .A2(new_n264_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n252_), .ZN(G1353gat));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n934_), .A2(new_n643_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n939_), .B1(new_n940_), .B2(new_n942_), .ZN(new_n943_));
  OAI211_X1 g742(.A(KEYINPUT126), .B(new_n941_), .C1(new_n934_), .C2(new_n643_), .ZN(new_n944_));
  XOR2_X1   g743(.A(KEYINPUT63), .B(G211gat), .Z(new_n945_));
  AOI22_X1  g744(.A1(new_n943_), .A2(new_n944_), .B1(new_n940_), .B2(new_n945_), .ZN(G1354gat));
  NOR2_X1   g745(.A1(new_n934_), .A2(new_n649_), .ZN(new_n947_));
  XOR2_X1   g746(.A(KEYINPUT127), .B(G218gat), .Z(new_n948_));
  NOR2_X1   g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n934_), .A2(new_n676_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n948_), .ZN(G1355gat));
endmodule


